MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       ~��@:��:��:��A��8��U��(�������U��G��X��7��:�����<����Ŷ�9��Rich:��        PE  L !@        � !  �        �     �                         �                              P� E   � �                            p �$                                                   �                           .text        �                   `.rdata  �-   �  0   �             @  @.data   ��   �  �   �             @  �.reloc  �?   p  @   P             @  B                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �D$V��L$W��N�:_ ���~�t�V�jRQ���Q_ ��t	W�&_ ��_��^� ��������������Q�_ YÐ�������H��t�T$�@jR+D$P�c_ � QV����^ ���D$tG�L$�T$jQR����^ ��u�NP�D$j h   P�R_ �D$^Y� �L$Q�^ �D$��^Y� ����A�A    Ð����V���H_ ���^Ð�Q�J_ YÐ���������8S�ك; VW�v  �L$H�j ��O�Q@P�Rh�������S  h`�jLj�~_ �����:  ���_ �����)  h'  ���6d Ph'  ���	d ����   h'  ���d Ph'  ����c ����   h'  ����c Ph'  ����c ����   h'  ����c Ph'  ���c ����   h'  ���c Ph'  ���c ��txj Vhb  j h�  ���` P�D$\�HQ�L$<�d Ph�  �T$(R���Wa �P�^ ��K��ۍL$���md �L$(�dd ���_ V�w^ ��_^��[��8� ���_ V�\^ ��_^2�[��8� ���������������	��u2�� �D$�PR��] H���@� ����������������	��t��] Ð����D$��0P�L$��k �L$ Qh���L$(�k P�T$R�ql P�| ���L$��k �L$ ��k �L$ �k ��0Ð���������D$��pP�L$$�ok h���L$�ak �L$tQ�L$�Sk �T$ R�D$P�L$Qh���L$p�6k P�T$`R��k ��P�D$LP��k ��P�L$8Q��k P�y{ ���L$0�-k �L$@�$k �L$P�k �L$`�k �L$ �	k �L$� k �L$ ��j ��pÐ���D$��0P�L$�j �L$ Qh���L$(�j P�T$R�Qk P�{{ ���L$�j �L$ �j �L$ �j ��0Ð���������D$��pP�L$$�Oj h���L$�Aj �L$tQ�L$�3j �T$ R�D$P�L$Qh���L$p�j P�T$`R��j ��P�D$LP�j ��P�L$8Q�j P��z ���L$0�j �L$@�j �L$P��i �L$`��i �L$ ��i �L$��i �L$ ��i ��pÐ���D$VQ�L$�$�n| �t$P���g jjj ����g ^Ð���L$�gf ��O�Q@P�Rh��j*h�  ���)] Ð��������L$�7f ��O�Q@P�Rh��j*h�  ����\ Ð��������L$�wf ��������L$��e ��O�Q@P�Rh��j h�  ���\ Ð���������V�t$W����e ��O�Q@P�Rh���΋��f �D$�D$Q�L$�$�b{ Ph�  �D$P����] ����y _^��Ð����V�t$W���`e ��O�Q@P�Rh���΋��e �D$�D$Q�L$�$�{ Ph�  �D$P���] ���y _^��Ð���L$�e ��O�Q@P�Rh��j h�  ����[ -b  ���@Ð��������������L$��HV��d ��O�Q@P�Rh����j�D$P�L$8�!_ Ph�  �L$$Q���_\ ����_ ���i �L$���g �L$�m_ �L$0�d_ ��^��HÐ�������������D$P�d YÐ�����V�L$�cz �D$(j �L$Q�T$R�L$�D$ �D$$    �D$(    �V{ �L$,P�L} �L$���q{ �L$�z �L$,������L$�dz ����^��Ð�������������O�T$�H@R�Qh�T$$���L$ QR�L$Q���D$    �D$    �D$    ��Z �D$�D$$�T$��L$�P�H���Ð���������������O�T$�H@R�Qh�L$��j Q���OZ �T$��Ð�����U������   �U��O�HTSV�uWRV�Q,��3���;�u	2�_^[��]á�O���   ���RT��;�u	2�_^[��]ÍL$4�x ��$�   P�Ή|$4�D$@   �|$D�|$L�|$H�|$P�|$X�D$\   �t$T�b ��$�   �L$@�Ή|$H�D$X   ��b ��O�M�D$<���   �PxP��$�   �e ��$�   �T$`�L$DR�Ή|$X��b ��L$4�P��O�T$8�|$L��T$0�L$0R���s{ ��t!��$�   �#e ��$�   ��\ 2�_^[��]��E�L$4�D$,    �D$(    �=��D$$    �D$p    �D$t    �D$x  �?�T$h�T$|ٔ$�   ٜ$�   �w �\$`�u�EN;ǉ|$��   �3��D$�|$�L$h�\$(�D$`�\$\�D$��O�T$\j �L$lj j R�\$4�H ��$�   P��$�   R�D$<Pj ��$�   SR�Q��P�@�L$@�D$@����(�T$�D$ F�z� �D$���F�h� �D$ ���F�V� ��EG;��|$�a����D$�M@;��D$�3������)z ��$�   �c ��$�   �[ _^�[��]Ð�������U������$��O�U�H@SVWR�Qh����j h�  ���bW �\$j hq  ���PW �\$j hs  ���>W �\$�X��D$�P�蕋 �\$$�D$�]�L$�C��D$�u�-H��   �D$� �=@�F;����\$�D$��|$�\$ ���D$�=8��\$�D$�=��\$��   �D$�L$�L� �L$�d$ �0�����t���D$(    �D$,    �%������Au���D$(    �D$,  �?��\$(�D$(�D$$��� �-��D$貊 �(�� �衉 �FG;��|$�h���_^�[��]Ð���������   ��O�HTS��$�   UVWjS�Q,��3���;�l$$�u  ��O���   ���PT��;��Z  �L$D�jt ��$�   Q�Ή|$D�D$P   �|$T�|$\�|$X�|$`�|$h�D$l   �t$d�o^ ��$�   �ΉT$P�|$X�D$h   �^ �D$L��O���   ���RxP��$�   ��` �L$l��$�   Q�ΉD$X�|$h��^ ���O�T$D�@�D$H�|$\��D$@P�͉T$D�Lw ��uwۄ$�   �L$D�D$0�D$,�=��D$(��$�   ��$�   Ǆ$�     �?�T$�T$t�T$x�\$|�s �\$l��$�   ����h����h�   Q�w �؃�;�u%��$�   �` ��$�   �IX _^]2�[�Ĵ   �;��k��|$��   �3��D$�|$�L$�\$,�D$l�\$�D$��O�L$j �L$ j jQ�\$8�B ��$�   R��$�   Q�L$<�T$@Rj Q��$�   R�P��P�@�D$d�D$d�T$`�D$`�L$\���D$\��(G;��h��|$�] |��D$@;ƉD$�V�����$�   O����   �   �L$�D$    ��L$������D1��   �֍��T$����֍��D$�L$��T$�"�D.������G��L$�����T$�$��`�葆 �`���*ЈG�� �T$��*Ȉ�L$�   �G�E�T$�U�;�� �L$|��l$�D$�@�D$H;Ɖl$�J���S�v �L$(���&u ��$�   �^ ��$�   �~V _^]�[�Ĵ   Ð��O�HT��  SU��$  VWjU�Q,��3���;�u_^]2�[��  Ë�O���   ���PT��;�u_^]2�[��  ÍL$|��p ��$�   Q�Ή|$|Ǆ$�      ��$�   ��$�   ��$�   ��$�   ��$�   Ǆ$�      ��$�   ��Z ��$�   �Ή�$�   ��$�   Ǆ$�      �[ ��$�   ��O���   ���RxP��$�   �>] ��$�   ��$�   Q�Ή�$�   ��$�   �
[ ���O�T$|�@��$�   ��$�   ��D$xP�ˉT$|�s ��t%��$�   �;] ��$�   ��T _^]2�[��  �ۄ$,  �L$|�D$\    �D$X    ݔ$�   �D$T    �=�ٔ$�   ٔ$�   ٜ$�   ��o ݜ$�   ��$0  ���D$0    �D$,    �D$(    �D$<    �D$8    �D$4    �D$$    �D$     �D$    �l  �$��( �D$  �?�L$�D$    �T$�D$    �D$�L$(�T$,�D$    �L$�D$    �T$�D$0�D$  ���D$�L$4�T$8�D$    �L$�D$  ���T$�D$<�D$    �D$�L$�T$ ��  �D$  ���L$�D$    �T$�D$    �D$�L$(�T$,�D$    �L$�D$    �T$�D$0�D$  �?�D$�L$4�T$8�D$    �L$�D$  ���T$�D$<�D$    �D$�L$�T$ �?  �D$    �L$�D$  �?�T$�D$    �D$�L$(�T$,�D$  �?�L$�D$    �T$�D$0�D$    �D$�L$4�T$8�D$    �L$�D$    �T$�D$<�D$  �?�D$�L$�T$ �  �D$    �L$�D$  ���T$�D$    �D$�L$(�T$,�D$  �?�L$�D$    �T$�D$0�D$    �D$�L$4�T$8�D$    �L$�D$    �T$�D$<�D$  ���D$�L$�T$ �  �D$    �L$�D$    �T$�D$  �?�D$�L$(�T$,�D$  �?�L$�D$    �T$�D$0�D$    �D$�L$4�T$8�D$    �L$�D$  ���T$�D$<�D$    �D$�L$�T$ �   �D$    �L$�D$    �T$�D$  ���D$�L$(�T$,�D$  ���L$�D$    �T$�D$0�D$    �D$�L$4�T$8�D$    �L$�D$  ���T$�D$<�D$    �D$�L$�T$ �D$$��$(  ��$,  N;�|$P�C  �3��D$P�|$@��ܴ$�   �%����L$�\$l�D$ ���\$p�D$$���\$t��݄$�   ٜ$�   �D$@��ܴ$�   �%��D$4��ٜ$�   �D$8��ٜ$�   �L$<ل$�   �D$(ٜ$�   �D$,؄$�   ٜ$�   �D$0ل$�   �D$l�\$Dل$�   �D$p�\$H�D$t�\$L�D$H�L$H�D$L�L$L���D$D�L$D�����������@t���D$    ����D$    �&�=��T$@�L$D�D$@�L$H�\$�D$@�L$L�\$����ٜ$�   �D$��ٜ$�   �D$��ٜ$�   �D$�����x��T$T�0�����t�D$T���\$T�D$��~ �p���O��$�   j �\$\�Q j j P��$�   Q��$�   P�L$lQj ��$4  SP�R��P�@��$�   ل$�   ����(�T$d�D$hF�S~ �D$d���F�A~ �D$h���F�/~ G;���|$@�����D$P@;ŉD$P��������m ��$�   �V ��$�   �`N _^]�[��  ÍI �" # �# A$ �$ c% �����������L$ �Ti �D$$�D$3�P�L$Q�T$R�L$�D$ �D$$�Nj �L$(P�Dl �L$�kj �L$ �i �L$(��L$ �ci ���Ð���������������L$ ��h �D$$�D$3�P�L$Q�T$R�L$�D$ �D$$��i �L$(P��k �L$��i �L$ �2i �D$(�L$ ���h ���Ð�������������� �L$ �th �D$(�D$3�P�L$Q�T$R�L$�D$$�D$(�ni �L$,P�dk �L$�i �L$ ��h ��P�@�L$�D$�D$�D$,����T$�T$�H�L$ �P�_h ��� Ð����������   VW��$�   ���ZS ����u_2�^�Đ   á�O�HpWV���   ����u��O�BpV�P����u_2�^�Đ   Ë�O�QHP�D$lP�RH��   �|$@�L$@Q�T$R�E  ��$�   �L$(�D$$�T$,��H�L$0�P�T$4�H�L$8�P�T$<�H�L$@�P �T$D�H$�L$���P(�T$�H0�L$_�@    �@    �@,    �P4�H8�@<  �?�^�Đ   Ð��SVW�|$W�0�����W�\$$�T���3���;މD$tl;�th���,R ��;�t[��O�HpWS���   ��;�u��O�BpS�P��;�t0��O�Q@P�Rh����Vh�  ���G ��thh��^�����_^2�[���h  Bh�  ���!G ��h  Bh�  ���\$�
G �D$ �|$_�p�p�p�p�p�p�p �p$�p0�p4�p<^�@(TI�?�@,  �?�@8II�[����D$�t$ ���X��؃�á�O�T$�H@R�Qh�L$P�D$PQ��  ��Ð�������������O�T$�H@R�Qh�L$P�D$PQ�  ��Ð�������������O�T$�H@R�Qh�L$P�D$PQ��  ��Ð������������D$�L$P��D Ð�D$��,S3�:�Vt�L$HSh'  �G U�L$$�D �l$@3�;�v2W�|$@�P�L$�Q �L$QV�L$0��G �L$��Q F��;�r�_��O���   ���   ;ÉD$D]u/��O���   �D$@P���   ���L$ �\$@�
D ^2�[��,ÍL$Q�L$�D$'  �\$�\$�te �T$@�L$DR�D$P��f �L$���e ;�t�L$ Qj���tG ��O���   �L$@Q���   ���L$ �\$@�C ^�[��,Ð������0V�D$ jP�0h ��jj
�L$(�F �t$\V�L$�P �L$Qj�L$(��F �L$�P V�L$�oP �T$Rj�L$(�F �L$�P �D$X��th)D �jj�L$(�F �D$@SQ�$j�L$,�&F �D$LQ�$j�L$,�F �D$TQ�$j	�L$,� F 3��D$�D$�D$P�L$P�D$'  �0d �L$d�� N  �T$R�L$H�t$�D$   �D$ �q �d �D$LP�L$(Q�L$t�T$LR�e ����ۍL$D���d �L$L�d ��[t�L$ �4B 2�^��0ÊD$d��t�D$8Q�L$p�$V�SE �L$ �
B �^��0Ð����@SV�D$4h�   P�f ��j j
�L$<��D �t$PV�L$(�O �L$$Qj�L$<�>E �L$$�%O V�L$(��N �T$$Rj�L$<�E �L$$�O h�   j�L$<�D �D$P�L$�D$'  �D$     �D$$    ��b �L$T�� N  �T$$R�L$�t$(�D$,�   �D$0�q ��b �D$P�L$8Q�L$d�T$R�Hd ����ۍL$����b �L$�b ��t�L$4��@ ^2�[��@ÊD$X��t&�D$LP�L$(�N �L$$Q�L$dV�DD �L$$�+N �L$4�@ ^�[��@Ð�����������<SV�D$0h�   P�Le ��3�Vj
�L$8�C h�   j�L$8�C jj�L$8�^C �L$Q�L$�D$'  �t$ �t$$��a �T$H�D$$�� N  P�L$�t$(�D$,�   �D$0�q �a �L$Q�L$P�T$4R�D$P�,c ����ۍL$���a �L$�a ��t�L$0��? ^2�[��<ËL$PV��? �L$0�? ^�[��<Ð���@SV�D$4jP�_d ��jj
�L$<�B �t$PV�L$(��L �L$$Qj�L$<��B �L$$��L V�L$(�L �T$$Rj�L$<��B �L$$�L h,D j�L$<�UB 3��D$�D$ �D$P�L$�D$'  �` �L$T�� N  �T$$R�L$�t$(�D$,   �D$0�q �y` �D$P�L$8Q�L$d�T$R�b ����ۍL$���` �L$�w` ��t�L$4�> ^2�[��@ÊD$X��t'�D$L� �L$`�\$$�@�\$(�@�D$$P�\$0V��A �L$4�j> ^�[��@Ð���\SV�D$4h�   P�c ��jj
�L$<�\A �t$lV�L$(�nK �L$$Qj�L$<�A �L$$�K V�L$(�KK �T$$Rj�L$<�{A �L$$�bK hD j�L$<�A 3��D$�D$ �D$P�L$�D$'  �R_ �L$p�� N  �T$$R�L$�t$(�D$,�   �D$0�q �&_ �D$P�L$8Q��$�   �T$R�` ����ۍL$���*_ �L$�!_ ��t�L$4�T= ^2�[��\ÊD$t��t9�D$hP�L$(�vJ �L$$Q�L$L�B �L$|PV�@ �L$H�TB �L$$�{J �L$4�= ^�[��\Ð�����������@SV�D$4h�   P�a ��jj
�L$<��? �t$LV�L$(��I �L$$Qj�L$<�.@ �L$$�J V�L$(��I �T$$Rj�L$<�@ �L$$��I hg j�L$<�? �D$P�L$�D$'  �D$     �D$$    ��] �L$P�� N  �T$$R�L$�t$(�D$,�   �D$0�q �] �D$P�L$8Q�L$`�T$R�8_ ����ۍL$���] �L$�] ��t�L$4��; ^2�[��@ÊD$T��t�L$\j V�5@ �L$4�; ^�[��@Ð�����`�L$h�A�I,�\$ �A(�I �\$h�D$ �d$h�A(�I�\$�A,�I�\$�D$�d$�\$�A �I�\$�A�I�\$�D$�d$�T$ �I$�D$�I�����I���0�����@��   �D$d��3��؉H�H��H�H�H�H �H�H�H,�H(�H$�L$$�T$$�L$(�L$,�ȉ�T$(�Q�T$,�Q�D$$  �?�L$$�H�D$(    �T$(�D$,    �L$,�P�H�D$$    �T$$�D$(  �?�L$(�P�D$,    �T$,�H�D$$    �L$$�H$�P �D$(    �T$(�D$,  �?�L$,�P(�H,��`��=�VW�A,�I�A(�I�A�I�\$ �A �I�\$�D$p�d$�	�����I���D$ �d$�I$�����\$8�A�I�\$�A�I�\$p�D$�d$�	�����I���D$�d$p�I$�����\$<���D$�d$�	�D$p�d$�I���D$�d$ �I�����\$@�����\$D�D$$���\$H�D$(���\$L�A$�I �D$l�A�t$8�I,�������\$P�A,�I�A$�I�����\$T�A�I�A �I�����\$X�A(�I�A$�I�����\$\�A$�I�A(�I�����\$`�A�I�A�I�   �����\$d���_^��`Ð���������������@SV�D$4jP�] ��jj
�L$<��; �t$PV�L$(��E �L$$Qj�L$<�!< �L$$�F V�L$(��E �T$$Rj�L$<��; �L$$��E jj�L$<�; 3��D$�D$ �D$P�L$�D$'  ��Y �L$T�� N  �T$$R�L$�t$(�D$,   �D$0�q �Y �D$P�L$8Q�L$d�T$R�4[ ����ۍL$���Y �L$�Y ��t�L$4��7 ^2�[��@ÊD$X��t'�D$L� �L$`�\$$�@�\$(�@�D$$P�\$0V�; �L$4�7 ^�[��@Ð�����L$j h'  �8 �L$��Ð�������D$�L$j  N  P�8 �L$��Ð����L$�D$ P�� N  Q�L$,�T$R�D$    �D$    �D$    �8 �D$�D$ �L$��T$�H�P�@  �?���Ð���8�L$ �; P�D$@ N  P�L$$Q�L$P��8 �L$ �< �T$@jh�   R�D$P�L$,�(< ���F �L$ �D �L$��; ���8Ð���������D$�L$ N  P�7 �����@Ð����D$�L$ N  P��6 �����@Ð����D$�L$ N  P��6 -�   ���@Ð��D$�L$ N  P�6 -�   ���@Ð���I��u:h��jh�   �VZ ����t���X  ����Iu� ��I    3�� j j j j�j�j j����H ������ �����������������0Vh'  �_ ��P�L$�B �L$�\C ��u�L$��B 3�^��0�h��j#j�Y ������t���\ ����3�h��L$�bB V�D$P����h��MB j �L$0Q�T$$R�D$HP��B ��Ph�q �Z ��$�L$$���KB �L$�BB �L$�9B ��^��0Ð�V���H\ �D$t	V�KY ����^� ����I��t�j���I    Ð����V����F �N��3 �N0�X�  �����^Ð�������������V���   �D$t	V��X ����^� ��V��N0����O�  �N�4 ����F ^Ð�������������j j h'  �K Ð��V��Wh�  �F   �F'  �F"'  �
H �Fj P�L$Q���D$'  �D$    �HH �Vj jh���h  ���R�D$P���D$ '  �D$$    �HH ��t��t�   �3��Nj jh���h  �Q�T$R���D$ '  �D$$    �	H ��t��t_�   ^���_3�^��Ð��������������D$������w�$��> �@   ø�   ø   ø   ø   Ð�> �> �> �> �> ���������� SUVW��~W�D$3�P�D$'  �\$�H ��u
_^][�� � �nU�L$Q���D$'  �\$��H ��u
_^][�� � �\$�^S�T$R���D$'  �H ��u
_^][�� � �D$4������	��   �$��@ hL�jAjT�V ����t����  ����u0h0��L$�0? �L$Q�O ���L$�J? _^]3�[�� � ��P�T$8�����M ��P��'  Q�]= �T$<P���R(��u?h��L$$��> �D$ P�7O ���L$ ��> ���$E �j���_^]3�[�� � j*W�N�u4 _^]�   [�� � ��~0��0P�(����M ��P��'  Q�W�? t΃�0���)D ��t���>R�������P�E -'  P�+�? t���0����C ��t���>Q������U ��P��'  R�|< P���W(_��^�]@[�� � �I J@ h@ p? ;@ �@ ;@ ;@ ;@ ;@ �@ �������������|$\  VW��uE�G��t>�w0���qC ��t0�GS�P�A����O��P��'  Q��; P���S(��[�_@^� _�   ^� ���SV��W�N0��C 3��^W���0 �����t#���C ��t�j���GW���c0 �����u݋���/ _^[ÐSVW�Y3�W���@0 �����t"����  ����t�WC GW���0 �����u�_^[� ��  ��t���B ��uօ�t�j���W���/ ���������V����V �N�$��
4 �N$�"#  2��FD�FF�FG�����^Ð������������V��N$�5#  �N�M4 ���V �D$t	V�S ����^� h��jjH�RS ����t���t���3�Ð���D$�D$     �L$ ����D$  �?�T$�D$    �L$�P�H��� ������8��OS�\$@VW��H@S�Qh���L$(���*3 Ph'  �T$R���h0 P�N�4 �L$�3 �L$(�}3 �FD�FE �P ���D$Hu�D$HP�P ��_^3�[��8� j P���vQ ��u�L$HQ�P ��_^3�[��8� �T$HR�pP ��_^�   [��8� ���������������V��L$�j j Q���FD�FE �FF�P���FF t�FG��u	�   ^� 3�^� �����t  SU��$�  ��V��W�FG��  ��$�  ����  ��O���   ���RP����O ���n  ��O�H@W�Qh�����L$<�|$(��1 Ph'  �T$`R���/ �L$<�92 �D$X�^P���3 ��t�L$XQ���*3 �FD�FE�FD���   jh�   ��$�   R�D$$P���,2 ���< �L$�: �L$Q��$�   �~$R���D$    �M!  ����  �FD�FF����  �D$����  �8 ��  �D$<P����1 Ph���L$|�w9 P�L$ Q�,: P�VJ ���L$�9 �L$t�9 �L$<�x9 �T$R�L$�:9 �D$P� J ���L$�T9 �T$�3�<(�D$ uB���3������I��v1�������Ѿ   I;�v�<)t���3�F�����I;�r���D$R�L$0��8 �D$����   hD��L$�8 �L$Q�L$0�9 �L$��8 �T$,R�I ����tojh�   ��$�  P�L$HQ���0 ���: �L$<�8 j NVj�T$HR�L$<�9 ���: P��$�  P��  ���L$<�U8 ��L$,Q�H ���L$,�=8 �L$X�0 _^]3�[��t  � �FF��u���
  �\$(3ҊVE3��FDSU�~$��RP�k!  ��t�3ɊNE3ҊVDSUQ��R�!  ��t���$�  �FD �FG �P�����$�  UP���V �L$X���|/ _��^][��t  � �������������V��L$j �RL � P�N$�7"  ^%�   � ����������������O��H  S��$P  UVW��H@S�Qh��$d  ��������   ��$d  j ��K � -'  tHtHuz�FD�FE�p�FD�FE �f�L$<�B. Ph'  �T$(R���+ �L$<�. jh�   �D$`P�L$Q�L$0��. ���8 �L$�6 �T$XjR���  ���L$ �e. ��$d  PUS����T _^][��H  � ���������O�T$�H@R�Qh���   � �����V�t$��Q�N�/ �   �FD�FE ^� ����������������A$Ð������������� Vh'  �R ��P�L$�5 hT��L$�5 j j �D$Ph�B j �L$(Qh�q �(R ���L$���5 �L$�5 ��^�� Ð����������D$��   S��$�   U3�V��$�   ��F�N�n�n�n�n �n$�n(�@��    WR�F�#L ��;ŉF(�O  P�FP����N��Q��K �V��R�F��K �F�F��P��K �NQ�F��K �VR�F$��K ���F��;ŉ~ ��  9n��  9n��  9n$��  ;���  �N����3��ʃ��N�~$����3��ʃ��F3�;���  �   �D$H�D$X�D$P�   �T$RQ�D$$�L$D�L$lP�L$DQS�D$0    �D$4    �D$L-   �D$T   �D$X'   �D$\   �D$d   �D$h   �D$l"   �D$t�   �l$|�dO����   9l$��   �F�T$ RPP�D$ PS�D$4�   �D$8�   �D$<s   �D$@z   �l$D�HO�N���V��;�tNP�LO�N���V��;�tSP�X��N���V9,�tZ�F �8�FG;������_��^][�Ĝ   � h���=�����_��^][�Ĝ   � h���!�����_��^][�Ĝ   � h��������_��^][�Ĝ   � h`��	�����_��^][�Ĝ   � �������SV��FW3�3�;�~\U�-ԑ�F ;�tE88t@�F��;�t6SP�ՋN��;�tP�ؑ�V���N��PR�PO�F��Q�TO�FG;�|�]�V$R�I �F P�^$�I �NQ�^ �I �VR�^�wI �FP�^�kI �N(�V��QR�^�ܑ�F(P�NI ��_�^(^[Ð���U����QSV��F�VW�}�~����QP�ԑhq  ����FPPj j ���h A  �đ�ȑh  ���̑h  �?j h  �?j h  �j �Б�F�D$    �P �L$Q���P��h�_ P�����D$�����h @�@j h  $@�\$�D$j h  �?j ���$�a! h   ���̑�v�N �F�V���v���D���$���F��$�����$�B���@�������\$���B���@�\$ �� �\$�@�\$�@�\$� �$��  _^[��]� ����������%������������V��F ��Wt_�|$�<8 tU�F$�<8 tL�N(��Rh�  ���h�  ����F��h�   Q�hOjh��  h�  ����V(��_^� _���^� ��������������V��F ��Wt7�|$�<8 t-�F$�<8 t$�N(��Rh�  ����F��h�   Q�lO_^� �����������0V��F ��W��   �F3�����   U�l$D�F�P �L$DQ���P��h�_ P�����F�P �L$Q���P��h�_ P������D$\����u�D$��t�   �3��N$�9�V �< t5�F$�<8 t,W�������L$@h P UQ�L$�}~  ���f����L$��  �FG;��U���]_^��0� ����������LV�t$T���q�  ����   �D$P�L$Q�T$R�D$`P���D$d    �D$    ��  ��uh�Ih����I�  ^��LÍL$Q��舍  h   �ȑ����T$R���ht�  ����D$TPj h  j����L$�T$Qh  ��    Pj���ht�  ������^��LÐ��������V��j�F �F    �D �F���F    �����^Ð���V���   �D$t	V��D ����^� ��V��FP����F ��D �����F    �	   ^Ð������V��N��t��P�F    ^Ð��������AÐ������������T$V��N�R�Pl��|�N��t��Pt��|�^� 2�^� V�������D$�L$�T$�F�D$�N�L$�V�T$�F0�N4�V@�����^� ��V���   �D$t	V��C ����^� �����������������   SUVW��Ǆ$�       �����L$d�D$4���  j jj �D$$P�L$$�D$t0��B  �L$��E  j�L$�D$���[G  Pj j �L$$�mF  �L$�Q�D$h��P�D���?I  �O�A��3�����   h��Vh��Vh��Vhl�VhT�Vh@�V�T$Dh0�R��H  ������4  P��H  ������4  P��H  ������4  P��H  �����4  P�H  �����4  P�H  �����4  P�H  �G�H��F;��[����O�A3���~3h��V�T$h�R�fH  �����\4  P�VH  �G�H��F;�|͍L$h��Q�9H  �W�B��3���~IhH�Vh�V�D$$h�P�H  �����4  P��G  ������3  P��G  �O�A��F;�|��T$h(�R��G  �G�H��3���~3h$�V�L$h�Q�G  �����3  P�G  �W�B��F;�|͍D$h��P�G  �O�A��3�����   Vhh�VhL�Vh0�Vh�Vh��V�T$@h��R�@G  �����63  P�0G  �����&3  P� G  �����3  P�G  �����3  P� G  ������2  P��F  ������2  �G�HF;��i����L$h��Q��F  �W�B��3����d  h��Vh��Vh��Vht�Vh`�Vht�V�D$DhX�P�F  �����x2  P�rF  �����h2  P�bF  �����X2  P�RF  �����H2  P�BF  �����82  P�2F  �����(2  P�"F  �G�H(�1������   �P$��h$�Ph�Vh��Vh��VhP�V�D$<h0�P��E  ������1  P��E  ������1  P�E  �����1  P�E  �����1  P�E  �����1  P�E  ��h$�V�L$h��Q�sE  �����i1  P�cE  �W�B��F;�������D$h��P�BE  �O�A��3���~3h$�V�T$h��R�E  �����1  P�E  �G�H��F;�|͍L$h��Q��D  �W�B��3�����   Vh��Vh��Vht�Vhd�VhX�V�D$@hH�P�D  �����0  P�D  �����0  P�D  �����0  P�D  �����v0  P�pD  �����f0  P�`D  �����V0  �O�AF;��i����T$h@�R�8D  �L$d����uS�D$8���tI�L$T��;�r���L$(�	�T$R+�PQ��$�   ��=  ��$�   P��$�   �.  j��$�   �   ��uM�L$4�9 tD�T$$��	�T$R�T$H�+��QP��$�   �=  ��$�   P��$�   �-  j��$�   �.�L$Q��$�   �F=  ��$�   R��$�   �-  j��$�   �<  ��$�   ��u�����H��؊��t
<�t�Ȉ�	Q�7= ����$�   U�wVj S�" ������   3�;�t	9] ��   ��W�R�P��}J�D$�H�D���D$\�D$��t�T$$�P��< ���D$\����L$�\$T�D$\��1  �   �D$�G�H�D���D$\�D$��t�T$$�P�< ���d$\��L$L;ˉ\$T�D$��t�
  ;�t�j����D$�H�D���L$d�D$d0���' _^]�[���   � �T$�B�D���L$�D$���;  �L$L�D$���r
  �L$�Q�D���L$d�D$d0��p' _^]2�[���   � �����@  V��F��u2�^��@  � ��$H  �D$DP�s�  ��u
^��@  � �V��$�   QR�T�������u
^��@  � �D$P�L$HQ��$�   R茍  �N��$�   PQ�+�������u
^��@  � ��$  R�D$P��$�   Q�P�  �T$R��$  P�.�  �N���jj�D$Pj �R4��}2�^��@  � �L$Q�T$HR�y�  �N���jj�T$Rj�P4��}2�^��@  � �D$P�L$HQ�Ĉ  �N���jj�D$Pj�R4����^��@  � �����������������  SUV��F��W�z  �F�~8Wh�  P藻�������]  �N�F9Ph�  Q�z��������@  �V�F:Ph�  R�]��������#  �F�n;Uh�  P�@��������  �N�F<Ph�  Q�#���������  �V�F=Ph�  R����������  �N��$�   PQ�j�������t.��$�   R��$�   P��  �N���jj��$�   Pj�R4�? �D$P    �D$T    �D$X    �D$\  �?��   �V�L$Qh4  R���������t>�N�D$Ph5  Q�O�������t$�D$�L$�\$P�D$ �L$�\$T�D$$�L$�\$X����~ Wj��h�  ����Rh�  ����F0�N4PQ��E �VPR��������t4�N4�F0Qh  h  PPjh�  �l ��N�Pj�RT�����N�j�D$TPj�R,�}  �D$`    �D$d    �D$h    �D$l  �?tX�V�L$Qh�  R��������t>�N�D$Ph�  Q�G�������t$�D$�L$�\$`�D$ �L$�\$d�D$$�L$�\$h�N�j�D$dPj�R,�F9���D$,    ��   �V�L$,Qh�  R��������t�F0�L$,�H��\$,�~$Wj��h�  ����Ph�  ����N0�V4�FQRP���������t,�N4�F0Qh  h  PPjh�  �! ��N�Pj�RT�N�j�D$0Pj�R�F:��Ǆ$�       Ǆ$�       Ǆ$�       Ǆ$�     �?�+  �V�L$Qh(
  R蝸������tG�N�D$Ph)
  Q��������t-�D$�L$ٜ$�   �D$ �L$ٜ$�   �D$$�L$ٜ$�   �n(Uj��h�  ����U Rh�  ���3�Ǆ$�   �  Ǆ$�   �  Ǆ$�   �  Ǆ$�   �  Ǆ$�   �  Ǆ$�   �  ��$�   �F0�N�+�S��P�F4PQ��������t"�F0�+V4Rh  h  ��PP�jP� C����|��E �N�Pj
�RT����N�j��$�   Pj	�R,�F<���D$@    �D$D    �D$H    �D$L    �  �V�L$Qh�  R裷��������   �~,Wj��h�  ����Ph�  ����N4�Vh   QR�E�������t4�F4Ph  h	  j h   h	  j h�  �����N�Pj�RT�L$���D$H�F=���щL$@�T$Dtd�V�L$Qh  R茶������tJ�N�D$Ph  Q��������t0�D$�L$�L$�\$@�D$ �L$�L$�\$D�D$$�L$�L$�\$H�N�j�D$DPj�R,�F�H3�ɿ   �4  3ۋ@�N�j�P��PG�R,�N�D$p    �D$t    �D$x    �D$|  �?�Q����$�   Qh�_ P�3�������tM�V�B���L$Qh�_ P��������t-ل$�   �L$�\$pل$�   �L$�\$tل$�   �L$�\$x�N�j�D$tP��PG�R,�V�D$0    �B�L$0Q��h�_ Q������D$<�����D$8  �?u�D$8    �F�D$4    �H�T$4R��h�_ R�����D$<����u�D$4���D$<    u�D$<  �?�N�D$    �Q�D$P��h�_ P�����D$� ��V�B�L$��Q��h�_ Q���@��=��\$,�����D$(� ��D$T�L$,�T$P����D$ j�D$ �L$(�NP�T$$���L$��P�\$4�G�R,�F�@�N�j�P��PG�R,�F�@�N�j�P��PG�R,�F�N�@��|$Gj�P�D$P�R,�F�HE��;�������N�A3ۅ�~&�N@S�,������t�N�)��PRG�UT�V�BC;�|�_^][��  � ��QV��L$�� �F��v	���sH�F�N3������L$H#��l ��^YÐ�������QV�1��t;�L$� �F��v	���sH�F�N3������L$H#��( ��t�j���^YÐ���������V��F��Wtb�F<���=ܑt�F,Pj�׊F:��t�N(Qj�׊F9��t�V$Rj�׊F8��t�F Pj�׋N�A3���~�N@W�����V�BG;�|�_^�V������3��F�F�F�P���^Ð��V���   �D$t	V�0 ����^� ��V��F��W�P�t3�F3���~#�F����t�j�R�F��    �FG;�|��F    �NQ�30 �F�����F    t=�F3���~!�V��P�0 �N����    �FG;�|ߋVR��/ ���F    �������_^Ð������������SU��E3�;�VW�E t7�E3�;�~�E��;�t�j�R�E���EG;�|�MQ�/ ���]9]�]t5�E3�;�~�U��P�f/ �M�����EG;�|�UR�L/ ���]�͉]�����t$(�D$$V�}WSP�0 �����M  ;�t9�A  ��E�P�R���.  �M�A��    R�E�. ����;��}�  �M������3��ʃ��9]~t�M��T$RS�P����   �t$��u������3������Q�). �M���U��������   ���3������+����������ȃ��EC;�|�3ۋM���    R�E��- ����;��}tX�M������3��ʃ��E3���~%�EVP�  �M���U������t�EF;�|�_^�E]�[��� �E _^]2�[��� ����V��F��Wu_2�^� �|$�D$WP�o�������u_^� �L$;N|�D$�T$�D$�NWR�QP�FRP������_^� ��SUV��F��Wu	_^]2�[� �F�l$ �\$3���~#�F���D$�UP�D$ PS�R��tˋFG;�|݄�t!�v��d}�� N  UV������F���N  |�_^]�[� ��������SVW���G��u_^2�[� �G3���~�\$�G���S���t܋GF;�|�_^�[� VW���G��t�G3���~�G����R�GF;�|�_^Ð������T$��'  |7�A��u2�� �� N  |#���N  �A��u2�� ���������P� �� ��������VW���G��t*�G3���~!S�\$U�l$�G���SU�R�GF;�|�][_^� ������VW���G��t�G3���~�G����R�GF;�|�_^Ð������D$U��j�E�?+ j(�E�5+ �L$�E�E�M�M���E �E    �E h��P�R����   �E�M�P�EP�R����   VW�L$Qh�����E�D$    �  ��t�|$��t�? u4�T$Rh�����  ��t�D$��t�8 u	�E��L$�U�:�|$��t�? u	����|$���3����Q�e* �|$����Ѓ�3��U���+����������ȃ��_^��]� ��]� ��������������V����   �D$t	V�k* ����^� ��S��U�l$�E�C3��C�C�M�K�UVW�S�C�h��}������Q��) ����ЉS�}3����+����������ȃ�j��) j(�C�) �S�C�M���A�B�I�J�u�{���
   �_^]��[� �����������V��FP�h��) �NQ�F    �) �VR�F    �~) ���F    ^Ð��� �����������Ð��������������2�Ð�������������D$�L$��VPQ�L$�y����D$��u�L$�h���3�^���j �( ������  �T$R���S  ������  �F����  �j���Pj�n( �����f  �L$Q����  �����P  �F����  �j���Rj(�2( �����*  �L$Q���  �����  �F���d  �j���Rj ��' ������   �L$Q���  ������   �F���(  �j���Rj$�' ������   �L$Q����  ������   �F����   �j���Rj0�~' ����tz�L$Q���  ����th�F����   �j���Rj,�J' ����tF�L$Q���  ����t4�F����   �j���Rj,�' ����t�L$Q���C  ����uh���3������L$����3�^��ÊF��u7�j���Rj��& ����t�L$Q���f  �L$���[�����^���3��L$�I�����^��Ð���$SV��F�H$W3���v>�\$4�N��D$P�FWP�R��|$�|$u�L$SQ��
 ����t�V�B$G;�r�_^2�[��$� �D$��T$8_^�
�[��$� ��������������$SV��F�H$W3���v>�\$4�N��D$P�FWP�R��|$�|$u�L$SQ�p
 ����t�V�B$G;�r�_^2�[��$� �D$8�L$_^��[��$� �����������������@$    � x�ËD$�T$P�A�IR�jPRh��� ������ �����������D$V��P�C����F�����t�F��t�   �F��^� 3��F��^� ������V���8   �D$t	V�[% ����^� ��V���� �D$t	V�;% ����^� ������u��������Q�D$��VW�|$���D$[��=tg�FWP���������t8�VW�L$QR���������u_^Y� �D$�^$����At�D$�^ ����t���D$��t���N�L$t�   �3��T$�F(�NWRP�F3ҊV,PQR���$���F$���\$���F �\$�D$@�$�=�����8_^Y� �����Ð�������������D$V��P������F����xu"�xu�H��u�H��u�H��u�   �3����F��   W�~ Wh�����������u�(kn΍~$Wh�����������u�(knN�~(Wh�����������u����=�L$Qh�����%�����_t�T$h��R�� ����u�   �3��N�VR�V�F,�R�P(��^� ��������V���   �D$t	V�;# ����^� ������u���������T$V��N�D$PQR��������t�N�j�T$R�VR�P^� �������������D$�T$P�AR�QjP�ARP�#������ ��������������D$S��P�C����K����C    �y�����Ct`�K�VW�D$P�CP�RP�KQ�i" �|$���3����Q��! �|$����Ѓ�3��S���+����������ȃ��_^��[� ��[� ���������������V���   �D$t	V��! ����^� ��V��FP�����! �����F    ����^Ð������������  SV��F��W��  ��$�  �D$P���D$  �?�D$    �D$    �D$    �D$     �D$$  �?�D$(    �D$,    �D$0    �D$4    �D$8  �?�D$<    �D$@    �D$D    �D$H    �D$L  �?��h  ��u_^[�Ā  � �F���|$tA��L$LQP�ϴ������u_^[�Ā  � ��$�   R�D$P�L$TQ�s  ����$�   �F��t=��T$LRP藵������u_^[�Ā  � ��$  P�L$PWQ��r  ����$  �F ��t��$�   RW�o  ����$�   �F��u��$L  PW�sn  ����$L  �N�F�jjWP�R4_^�[�Ā  � �����������D$SV��P�����N2��ؔ�^�Qh��R�& ����u��F�F�^�^�^�^ ��^[� �F�Hh��Q�� ����u��F�F �F�^�^�^��^[� �V�Bh��P�� ����u��F�F�F�^�^�^ ��^[� �N�Qh��R� ����u��F�F�F �F�^�^��^[� �F�Hh��Q�Z ����u��F�F�^�^�^�^ ��^[� �V�Bh��P�' ����u��F�F �F�^�^�^��^[� �N�Qh��R�� ����u��F�F�F�^�^�^ ��^[� �F�Hh��Q�� ����u��F�F�F �F�^�^��^[� �V�Bh��P� ����u��F�F�F�^�^�^ ��^[� �N�Qh��R�[ ����u��F�F�F �F�^�^��^[� �F�Hh��Q�( ����u��F�F�F�F�^�^ ��^[� �V�Bh��P�� ����u��F�F�F�F �F�^��^[� �N�Qh��R�� ����u��F�F�^�^�^�^ ��^[� �F�Hht�Q� ����u��F�F �F�^�^�^��^[� �V�Bhh�P�\ ����u��F�F�F�^�^�^ ��^[� �N�QhX�R�) ����u��F�F�F �F�^�^��^[� �F�HhD�Q��  ����u��F�F�F�F�^�^ ��^[� �V�Bh,�P��  ����u��F�F�F�F �F�^��^[� �N�Qh�R�  ����u��F�F�F�F�F�^ ��^[� �F�Hh��Q�]  ����u��F�F�F�F�F �F��^[� �����������V���   �D$t	V�� ����^� ���ؔ�����������  SV��F��W�N  �F����$�  �D$  �?�D$    �D$    �D$    �D$    �D$   �?�D$$    �D$(    �D$,    �D$0    �D$4  �?�D$8    �D$<    �D$@    �D$D    �D$H  �?�|$t7�D$LPS����������   ��$�   Q�T$R�D$TP�+m  ����$�   �F��t/�L$LQS迯������tl��$  R�D$PWP��l  ����$  �F ��t��$�   QW�Fi  ����$�   �F��u��$L  RW�h  ����$L  �N�V�jjWR�P4_^[�Ā  � ���D$��VW�|$(���D$[��=�D$[��=�D$[��=�D$[��=��   �FWP����������   �VW�L$QR��������u_^��� �D$�������uw�D$�������Atf�D$�������uU�D$�������AtD�D$�������u3�D$�������At"�D$�������u�D$�������Au���D$ ��t)���N��T$�Q�T$�Q�I�T$�L$t�   �3��T$$�NWRP�FPQ�T$R辴����_^��� ����D$��VW��P�����N����yh�W�� ����t:h�W�� ����t(h�W��� ����th��W��� ����t3���   ���F�   t�V9Ju�   �3����Ft!�T$R�V�L$�NR�V�D$    �R�P0_��^��� ���V���   �D$t	V�+ ����^� ������e���������D$��   ��S��$  VW��|$tP�FSP��������t"�VS�L$QR�B�������u_^[��   � ����$  ��t���~$t�   �3���$  �VSQP�FRPW舴����_^[��   � ����������D$U��P�����M�E ��E$    �I��t��t	��t3���   ���E��   �T$R�Mh,����D$    ������t�D$��u%�D$Ph$���������t�D$��u�D$�I�M$VWQ�� �|$���3����Q�a �|$����Ѓ�3��U$���+����������ȃ��_^��]� ��]� ����������V���   �D$t	V�k ����^� ��V��F$P���N �����F$    ����^Ð������������4  SUV��W�k Uj����K��$L  �D$DPQR�r���������  ���3��|$D��эD$DI��t	����  �t@�T����:u��t�P��:Vu������u�3��������t�D$DPhD��ӓ����_^][��4  � �L$ ��i  j���̍T$+R�D$\P�  �L$4�;j  ��u�L$DQh4�舓�����8  �D$)��t�U Rh�  ����L$ �s  �  �D$*��t�E Pho�  ����L$ �s  ��   �t$0�F���D$u�L$ �Mp  ��   �D$�\$���8����\$<�8����D$���t$<� ���$ �D$�D$��% �\$����@t]�F�\$�8����D$���t$<� ��$ �D$�D$�% �\$����@t!�M Qh�  ���h�  j �L$(��p  ��U Rh��  ����L$ �Xr  �U �K�R�SR�PT�L$ �h  _^][��4  � ���� Qj�ܑÐ���D$�T$P�ARP荮����� ��������D$V��P�S����N�0��y����V��^� �������V���   �D$t	V�{ ����^� ���0������������VW�|$��N�D$P3ҊV3��FQ��RP�\  ��uh�Ih\����[  _2�^��� �N�j�D$P�FP�R,3Ʌ���_��^��� �������D$��VW�|$��t"�FWP���������t�D$��t�   �3��L$�VWQP�FRP������_^� �D$V��P�3����N�L��Qh��R�� ��������Fu�F�Hh��Q�� ����u�V�zu�   �3����FtF�D$Ph�����D$    ������t$�L$h��Q�Q� ����u�   �F��^� 3��F��^� �V���   �D$t	V�� ����^� ���L�������������D$��VW�|$(���D$[��=�D$[��=�D$[��=�D$[��=tF�FWP胶������u���D$ ��t)���N��T$�Q�T$�Q�I�T$�L$t�   �3��T$$�NWRP�FPQ�T$R謳����_^��� ��D$��VW��P�����N�l��yh�W�8� ����t=h�W�&� ����t+h�W�� ����th��W�� ����t�   �3����F�   t�V9Ju�   �3����Ft!�T$R�V�L$�NR�V�D$    �R�P0_��^��� ���V���   �D$t	V�K ����^� ���l�����������T$��V��N�D$PQR�W�������t�N�j�T$R�VR�P,^��� ������SUV�t$���W3���{�{�{�N�����;�s��;�u`;��v��� ����  �C+�;�s��;�v/�K�+�P�1RQ��" �k��W+�U���/  ��tU���  ���  _^]��[� ;�vK;�uG�F;�u����x��s5�{�{�{�F;�u����C�N�K�V�S�H�_^���H�]��[� jU���  ��t'�v;�u����{�͋����ȃ��U���o  _^]��[� �������D$SU��V3��M W�|$3�����u�u�u���I�ك��v�� �M;�t%�A���t<�t;�uA�ȈA�V���)  _^��][� ;�uj���  _^��][� �E��w;�sj����  S���=  �}�t$�ˋ����ʃ��E_�]� ^��][� ���U��j�h �d�    Pd�%    ��   SVW�e���8���3�3��}��  :��H  ��@Ƌ@ �Eԋ��  �M���� ��W�j  jP�M��� ��;�uD�M��I� ����  �=�I;�u*j� ��;�t
S���	  �3�P�/4  ����I���M��,� �M�;�t����;�t�j�����H�L1��   �M؉]�;�u3���HΉ�x����P�2�P0�U��@(�E��]̋Ủ�|����E���]S�]�SQP�E�P�M�Q���R�EĄ�t:�E�   �1��8�����JȋA���Q(��u��jP��� ��� Ë�8����E������}��J΅�t�AǋQ(��u��j P�� �� ��uL��H�1�@t>3��@u�@(����R,���u�   ��H΅�t�AǋQ(��u��j P�A� �ƋM�d�    _^[��]� �E����E�P�M��" �E�,�h���M�Q�J' �����,���" �������Q�L$�" h���D$P�D$,��' ������������V���,��" �D$t	V�u ����^� �������������D$V��P�A" �,���^� �������QV��L$�v� �> u��W@��W��6�L$��� ��^YÐQV��L$�F� �F���s@�F�L$��� ^YÐ����������2�Ð�������������Ð������������QV����q4��t;�L$��� �F��v	���sH�F�N3������L$H#��a� ��t�j���^YÐ������ ����������3�Ð���������������Ð�����������V���P���u�^ËF,��v��H3҉�^��Ð�������QSUVW�|$3����ىD$~z�l$�C�0��tG�K,���~>;�}�ǋȋ������ʃ��L$�|$ȉL$�K,)�K�+��Љ|$������P���t�L$�E EAO�L$�|$����D$_^][Y� ���������QSUV�t$3���W�ىD$~�l$�C �8��tI�K0���~@;�}�Ƌȋ������ʃ��L$�|$ȉL$�K0)�K �+��Љ|$����!�3ɊM Q���P���t�L$EAN�L$�t$����D$_^][Y� ����V�t$��������F���N�L$��� �XX�L$�V�x� ��^� ���V�t$��������F���N�L$�� �XX�L$�V�8� ��^�  ������ ������������D$�����UVW��u_^3�]��� �M �	��t&�U0�2�<;�sN�2�m �M _�Q�U ^�]��� �EDt_^���]��� �E�8 u3��|$��U0�u�>�+���D$���u@��t$��y3�SP�I ������v!�E�0�ϋ������ʃ��t$�|$��M@�   ;�~�E@�EDt�E�Q�_ ���MD�����MDu#�U�]<��E ��M0�1�U��E��M,�9�r�E�8�M<��+�ʋU�M<��E � +���+�:�M Ë�+Љ�E0։�EDt�M��U��E,�     �"�U�E� �:�M �	+�É�U+ȉ�E,A��E0��m �M �D$[_�Q�U ^�]��� ����������A� ��Vt@�Q;v9�T$���t:P�t�ADu%�A,� �A�0N����0t�A�^���� ^3�� ^���� ���������������SV�q���WtO�y,����;�s
3Ɋ_^[����ADu2�Q ���t);�w9A<v 9Q<s�Q<��A<+3��A�_3��^[�_^���[Ð��������������Q ���SVWt9A<s�A<�\$����   �A�0����   �D$��u�Q�:�A<�T$+���+��u����   �Q�:�T$��+�������   �T$����   �A� �y<+�;���   +Ƌq,�>�+��>�q�>����>��   �y �����   �A�0�A0� É7�I0+Ɖ�m��te�2��t_�D$��u�Q��A<�T$+�����u�Q��T$��+�����u*�T$��|"�A� �y<+�;�+Ƌq0�>�+��>�I �����t$����N���L$�V�� �XX�L$�F�/� _��^[� ���������D$�T$SVW�y Ћ��t9A<s�A<�����   �\$,��tV�A�0��tM��|z�A� �y<+�;�l+Ƌq,�>�+��>�q�>����>tT�y ���tK�A�0�A0� É7�I0+Ɖ�4��t,�?��t&��|"�A� �q<+�;��q0+ǋ>�+��>�I �����t$����N���L$,�V�� �XX�L$,�F�3� _��^[�  ������������V�q���P�N�D
����0��� �D$t	V� ����^� �����������V���0��� �D$t	V�� ����^� ������������QVW������w4��t;�L$��� �F��v	���sH�F�N3������L$H#��n� ��t�j����D$t	W�v ����_^Y� �����������VW�y���H�wP�D1����F��F���t�V��P�3 ���f���N��F�    �F��������N��Q�D2������0��� �D$t	W�� ����_^� ����QV���FD���t�F�Q�� ���ND���W�F<    �ND����~4��t;�L$��� �G��v	���sH�G�O3҅��L$J#��T� ��t�j����D$_t	V�[ ����^Y� ��D$��V��t#�F��t�H����t
<�t�Ȉ�	Q�% ���F    �F    �F    ^� ���������Q�D$��VW���D$    t����G(    �G0���H�D$���9��tI��r�D$��ΉF(�F,    �F0 �� �F(��u�F��j ��P���� �D$��t���� ��_^Y� ��V���FDt�F�Q�\  ���FD����F<    �FD^Ð���������L$�3Ɉ�H�H�H� ���������D$S�\$U��V3�����M �u�u�uv��� �M;�t$�A���t<�t;�u?�ȈA�V������^��][� ;�uj���q���^��][� �E��w;�sj���T���S���  �t$W�}�ˋ����ʃ��E_�]� ^��][� ��D$�A�I� � ���������������SVW�|$�����v�1� �F3�;�t*�H�:�t#���t;���   �ɈH�_�^�^�^^2�[� ;��L$uU:�t@;�t+�H��:�t<�t�Ȉ_�^�^�^^2�[� Q���  ��_�^�^�^^2�[� ;�t�^�_^2�[� :�t\�N��w;�s];�t3�H��:�t!<�t�ȈW�Ή^�^�^�w  _^�[� Q�i�  ��W�Ή^�^�^�U  _^�[� 9~sW���@  _^�[� ��������S�ً�H��H��VWuO�p,��tH��B�L0�3���u�@(����R,���u�   ��H΅�t�A�Q(ǅ�u��j P��� ��Q�L_3���^��[Ð����������VW���� �L$�F4��� �=�W�L$��� �G���s@�G�L$�S� �L$�J� �F�F�N�N�V�V ����F�F�N$�N,�V(�V0�     �F �     �N0�    �V�    �F�     �N,_���    ^��Ð������D$S��3�U�l$;�K8�K<�C@    �CD��   ��<��   ;��}3�VWP�_�  �t$�͋������ʃ��(���K<�CD_^u�S��K��S,�*�CDu*�K��S ��K0�)�S�: u�K��S��C,�     �CD��]�CD[� �S�
�C��S,�
�C��S �
�C0]�[� ���������L$3���u�   ��u��� �����U��j�h0�d�    Pd�%    ��@SVW�e��ى]��E�����u���v�E���E�    �F�E؅�}3��E�P�I�  ���E��'�E�E����}3�P�,�  ���E踰� Ë]��u��E������C��v";�v�Ƌȋs�E�x�����ʃ��u�{�C��t�H����t
<�t�Ȉ�	Q�'�  ���C    �E�@�C�@� �s;�w���s�K�1 �M�d�    _^[��]� ������������SU��M3�;�VW��   �A�����   <���   �ȈA�����3����U�U�U���I�ك��v�� 3ҋM;�t!�A���t<�t;�u9�ȈA�R������_^][�;�uj������_^][ËE��w;�sj�������S���9����}�ˋ����ȃ��M�]� _^][Ð������U��j�h@�d�    Pd�%    ��   SVW�e�3҉U�}���3����I���}܋u��H�D1;�~;�v+ǉE���U��������މ]��u
�   �  �E�    ��B�D0�E�%�  ��@��   �E���vp��Q�2�P0�U��H(�M��U��A � �E���t,�E��y0��;�s�H��I ��E��x�9��E�%�   ���E�%�   P�R�E��E��������u8�M��E����   �}܋�Q�L2(�M��W�UR�P�E�;�t�E�   ��M��M����E���vp��H�1�P0�U��H(�M��U��A � �E���t,�E��y0��;�s�H��I ��E��x�9��E�%�   ���E�%�   P�R�E��E��������u#�M���AƉ�x����P��|����@    �3�M��b����E��IȋA���Q(��u��jP�9� �-� Ëu�E������]�U��H΅�t�AQ(��u��j P�� �
� ��uL��Q��@t>3��@u�@(����R,���u�   ��H˅�t�AǋQ(��u��j P�� �ƋM�d�    _^[��]Ð���������D$��@V��h��L$�F���� �L$�U� ��^��@� ���������������,U�l$@V�E P�L$�  �L$�D� ��W����jP�L$�M� ����uE�L$�� ���2  �5�I��u*j�c�  ����t
V���  �3�P��  ����I���L$�v� �L$��t�������t�j����D$LSWj �L$0�D$0�����E��@uV�\$T����T$4����+ʃ�0��w�3� �T$4�rj V�L$4�������t~�L$0�T$4���V�L$0��������a�D$T��t+��D$P���R���Qj �T$$R�L$8��  j�L$ �)��L$Q���P���Rj �D$$P�L$8�  j�L$ �Z����E���\$4~
;�v+Ë��3��M�l$P���  ��@t1���T$D�D$H�T$�D$vU�L$�  Ou�\$4�L$�D$3���D$H�L$D�t$0��u����ۉL$D�D$Hv3ɊQ�L$H��  FKu���T$L�D$D�t$H�B    �D$v��tU����  ���u�D$Ou�|$@�L$��L$0�ɉwt&�A���t<�t�ȈA���_[^]��,� IQ��  ����_[^]��,� h���L$�   h���T$R�� �����V�D$��P�$ �,���^� ��������D$V�0W���L$�7�� �F���s@�F�L$�� ��_^� ���������������SUV�t$W�|$9w��s�� �G�L$��+�;�s��;���   �E�=���;�s��� ��������E+�;�s����v6�M�+�P�9RQ� �u��j +�V���Q�����t
�E�u� �t$�͋������E;�s�����K  �M+�P�9RQ�� �u��j +�V���������!  V�������_^��][� 3�;�vp;�ul�G;�u����x��sZ�E;�t�H����t
<�t�Ȉ�Q���  ��3҉U�U�U�G;�u����E�O�M�W�U�H�_��^�H���][� ���]  ;�s�� �M��t%�A���t<�t��uA�ȈA�S���A���_^��][� ��uj���+���_^��][� �E��w;�sj������S���U����G��u����}��ˋ����ȃ��M�]� _^��][� ��A V�0��t*�A0�W�<2;�_sJ��A ��Q��D$�%�   ^� �T$����   R�P^� ����������|SV��$�   �N�� W�D$$%�D$%t	�D$%+�D$&��t� #@��� l��   @��   u�o���   t�d��р�������@ ��$�   P�L$(Q�T$PR�B ��$�   ����$�   �D$8�D$T��<+�|$�\$H�L$0t(<-t$<0u�D$I<xt<Xu
�D$   ��D$    ��D$   �� V�L$�����L$ �&� ��W����jP�L$�/� ����uE�L$�v� ����  �5�I��u*j�E�  ����t
V���v  �3�P�  ����I��U�L$$�W� �L$�����T$<R���s  ����P�l$@��D$$���t�ŀ8 �����D$tj��u����E <���D$ tS��~O�T$����+�;�s@�T$+�+�BR�|4P�D4QWP�X �L$ ���,�EA���L$~E�E <�|$�D$u���$�   �A��~;�v+ǉD$��D$    �A%�  ��@��   =   t$�L$��$�   ��$�   Q��$�   RPQ�T$,R�J�L$�D$��$�   Q��$�   R��$�   P+��\X�D$XPQR�D$4P�|$0��  �H���QR�D$,P�D  ��P���L$0�T$4�D$    �D$��u#�D$4�L$0WSPQ�T$@R�~  �0�x���   h�S�
 �L$8��D$<USPQ�T$HR�N  �0�x�D$0���+ŉD$tZ�D$$��t�D$$jPW�L$(VQ�  �0�x��Ch�S�)
 ��USW�T$DVR��  �0�x�L$0���+Ń��ȉL$u��T$��$�   ��$�   RPWV��$�   V�A    �D  ��j�L$@�����]_��^[��|� h���L$0�|���h���L$0Q�c	 ���������������|SV��$�   �N�� W�D$$%�D$%t	�D$%+�D$&��t� #@��� l��   @��   u�o���   t�u��р�������@ ��$�   P�L$(Q�T$PR�R	 ��$�   ����$�   �D$8�D$T��<+�|$�\$H�L$0t(<-t$<0u�D$I<xt<Xu
�D$   ��D$    ��D$   �� V�L$�����L$ �6� ��W����jP�L$�?� ����uE�L$�� ����  �5�I��u*j�U�  ����t
V���  �3�P�  ����I��U�L$$�g� �L$������T$<R���  ����P�l$@��D$$���t�ŀ8 �����D$tj��u����E <���D$ tS��~O�T$����+�;�s@�T$+�+�BR�|4P�D4QWP�h�  �L$ ���,�EA���L$~E�E <�|$�D$u���$�   �A��~;�v+ǉD$��D$    �A%�  ��@��   =   t$�L$��$�   ��$�   Q��$�   RPQ�T$,R�J�L$�D$��$�   Q��$�   R��$�   P+��\X�D$XPQR�D$4P�|$0��
  �H���QR�D$,P�T  ��P���L$0�T$4�D$    �D$��u#�D$4�L$0WSPQ�T$@R�
  �0�x���   h�S� �L$8��D$<USPQ�T$HR�^
  �0�x�D$0���+ŉD$tZ�D$$��t�D$$jPW�L$(VQ�
  �0�x��Ch�S�9 ��USW�T$DVR�	
  �0�x�L$0���+Ń��ȉL$u��T$��$�   ��$�   RPWV��$�   V�A    �T
  ��j�L$@�����]_��^[��|� h���L$0����h���L$0Q�s ��������������D$��lSUV�p��W�H�� u�   ��$�$   ���H�� �D$ %�D$!t	�D$!+�D$"��t� #@� .@� *�� 0  @��    u�f���   ��I�����g���$�   �@ ��$�   PQW�T$,R�D$@P�@ ��$�   +���$�   �؋B�΋�$�   ������$�   �L$�l$0~�;�v
+�+ÉD$���$�   �D$    �D$��$�   �I���  ��@��   ��   t6����$�   �t$�T$v����$�   P�L$�c	  Nu�t$�|$�   ��vN�L$0��+t��-u@��$�   Q��$�   ��$�   ��$�   �	  ��$�   ��$�   �D$K�l$1��$�   ����$�   ��$�   v����$�   P��$�   ��  Nu鋴$�   ��$�   �D$    S�� ��RU�> �؃�����   ��$�   �� P��$�   �z���j��$�   j Q��  ��$�   ���ɉD$t������t�j���+�C�C�PUW�L$4VQ�"  �L$,�0��x���Rj��$�   ��$�   PW�L$4VQ�  �0�x��$�   ���+É�$�   ��$�   RjeU�z ������   +�@�؋D$Pj0�K�QUW��$�   VR�  �H���QR��$�   P�  ��$�   �Q�����D$    ��u���P� jQRP��$�   Q�M  �0�x��$�   ���+É�$�   �T$��$�   Rj0PUW��$�   VQ�  �P� ��RP��$�   Q�  ��$�   �Ћ�J��$�   �B    �T$$R��$�   RQPV�\  ��(_��^][��l� ��������������D$��lSUV�p��W�H�� u�   ��$�$   ���H�� �D$ %�D$!t	�D$!+�D$"��t� #@� .@� *@� L�� 0  @��    u�f���   ��I�����g���$�   �@ ��$�   PQW�T$,R�D$@P�l ��$�   +���$�   �؋B�΋�$�   ������$�   �L$�l$0~�;�v
+�+ÉD$���$�   �D$    �D$��$�   �I���  ��@��   ��   t6����$�   �t$�T$v����$�   P�L$�  Nu�t$�|$�   ��vN�L$0��+t��-u@��$�   Q��$�   ��$�   ��$�   �K  ��$�   ��$�   �D$K�l$1��$�   ����$�   ��$�   v����$�   P��$�   �  Nu鋴$�   ��$�   �D$    S� ��RU�j  �؃�����   ��$�   �� P��$�   ����j��$�   j Q�%  ��$�   ���ɉD$t������t�j���+�C�C�PUW�L$4VQ�N  �L$,�0��x���Rj��$�   ��$�   PW�L$4VQ�  �0�x��$�   ���+É�$�   ��$�   RjeU��  ������   +�@�؋D$Pj0�K�QUW��$�   VR��  �H���QR��$�   P�D  ��$�   �Q�����D$    ��u���P� jQRP��$�   Q�y  �0�x��$�   ���+É�$�   �T$��$�   Rj0PUW��$�   VQ�@  �P� ��RP��$�   Q�  ��$�   �Ћ�J��$�   �B    �T$$R��$�   RQPV�  ��(_��^][��l� ����������D$��TSVWP�L$ h�Q�$�  �T$|�؋B����~
;�~+Ë��3ɋR���  ��@�L$xUtp�ɋD$l�t$p�D$vT����tF�N ���t&�F0��,;�sI��F ��Q��D$x�%�   ��L$x����   Q���P���u�D$Ou��D$3ɉL$|��t$p�D$l�ۍ|$ �D$vi�\$��tL�V �����\$lt&�N0��,;�sJ��F ��Q��D$l�%�   ��L$l����   Q���P���u�D$�D$GH�D$u��L$|�ɋT$t�D$�B    �D$l]vT����tF�N ���t&�F0��;�sI��F ��Q��D$t�%�   ��L$t����   Q���P���u�D$hOu��D$d�T$h_��p^[��T� ���������D$V����t	V�z�  ����^� �Q�D$��V�t$voSUW�|$$�D$��tL�F � ����\$(t&�N0��,;�sJ��F ��Q��D$(�%�   ��L$(����   Q���P���u�D$�D$GH�D$u�_][�D$�T$��p^YÐ���D$��V�t$vZS�\$UW����tB�F ���t$�F0��,;�sI��F ��Q��È%�   ���ˁ��   Q���P���u�D$Ou�_][�D$�T$��p^Ð��������������Ð���������W���O��tG�A V�0��t(�A0�S�2;�[sJ��I ��B��D$�%�   ��D$�%�   P�R���^u���_� �������V�t$V�P��^� �����������������TVW�L$�� �L$��� �5�W��u�5�WF�5�W�5�W�L$�r� �|$`jV����� �����9  �D$h���>  ��� � ���/  �5�I���  j���  ��������   SUh��L$(�F    ���� ��  ���V�H��V�X���3������I��GW��  ������v
��M ECOu�����F3�� ������I��GW�e�  ������v��+ˊ�COu�j h��n��  ���L$$�F�� ][�3��L$`��� �L$h�5�I�� �F���s@�F�L$h�=� h� ��  ���L$`�'� �5�I�L$�� _��^��TÍD$hP�L$�D$l�����  h���L$Q�D$,��z�  �����AÐ������������AÐ�����������Q�I�D$SU�l$V3��L$W������E 3��u�u�u���I�ك��v�� �M;�t&�A���t<�t;�uC�ȈA�V���3���_^��][Y� ;�uj������_^��][Y� �E��w;�sj�������S���E����}�t$�ˋ����ʃ��E_�]� ^��][Y� ����������Q�I�D$SU�l$V3��L$W������E 3��u�u�u���I�ك��v��� �M;�t&�A���t<�t;�uC�ȈA�V���c���_^��][Y� ;�uj���L���_^��][Y� �E��w;�sj���-���S���u����}�t$�ˋ����ʃ��E_�]� ^��][Y� ����������Q�I�D$SU�l$V3��L$W������E 3��u�u�u���I�ك��v��� �M;�t&�A���t<�t;�uC�ȈA�V������_^��][Y� ;�uj���|���_^��][Y� �E��w;�sj���]���S�������}�t$�ˋ����ʃ��E_�]� ^��][Y� ����������V��FP���^�  �NQ�U�  �VR�L�  �D$�����t	V�5�  ����^� �������������D$��@SUV��Wh��L$�C���b� ���  ���S�H��S�h���3������I��FV�p�  ������v
�M �GENu�����C3�� ������I��FV�@�  ����v��+��U �/ENu�����C3��������I��FV��  ������v��+͊E �)ENu��L$�{�j� _^]��[��@� ���������������QV�L$�h� �t$�L$�5�I�U� �F���s@�F�L$��� h�� �\�  ���L$��� ��^YÐ�QV�L$�� �t$�L$�5�I�� �F���s@�F�L$�� h� ��  ���L$�v� ��^YÐ���V�L$��� �5�I�L$�� �F��v	���sH�F�N3������L$H#��-� ��t�j����L$��I    �� ^��Ð�����������V�L$�V� �5�I�L$�G� �F��v	���sH�F�N3������L$H#��� ��t�j����L$��I    �� ^��Ð���������S�\$V���W3������I��FV�4�  ��������v	��ACNu���_^[Ð����������TXS���u
âTX�8   �UX��u
âUX�3   �VX��u
âVX�.   [Ð�����������h@� ��  YÐ���h@� �o�  YÐ���h@� �_�  YÐ���Ð���������������D$S3�V���^�^�^�^�^�^ �^$�^(�^,�d  �NhD���jQ�q�  ��;ÉF��   �VS��RP���  �FhD���jP�B�  ��;ÉF��   �NhD���jQ�!�  ��;ÉF��   �VhD���j R� �  ��;ÉF��   �FhD���j$P���  ��;ÉFtc�NhD���j(Q���  ��;ÉF tF�VhD���j,R��  ��;ÉF$t)�Nj���QP�,�  �VhD�j1R�|�  ��;ÉF(uh(��xS������^[� �NSQP���  �����)  �F,��^[� ��������������V��F(W3�;�t	P�M�  ���F$;ǉ~(t	P�:�  ���F ;ǉ~$t	P�'�  ���F;ǉ~ t	P��  ���F;ǉ~t	P��  ���F;ǉ~t	P���  ���F;ǉ~t	P���  ���F;ǉ~t	P���  ���~_^Ð����������������O���   V�t$���R4��uB��O���   ���R(��u.��O���   ���R0����t��O���   ���R(��u��3�^� ���  SU��M �E    �E    谹  �؅���  VW��O���   ���R=�  ��  ��O�HHj hIr S�Qx�����D$tH��O�J@P�Qh����j h�  ���
�  j ��h�  ���D$#���  ���D$�D$���g  �E���N  �U����O�HH��$   SR�QH���E���   ��$�   �ل$�   �MS��U�Eل$�   ���\�M�Uل$�   ���\�E�M���D  �?��O�BH��$l  Q�PH��   �|$P��D$t�L$t�D$x�L$x���D$|�L$|�������������@t���D$$    ����D$     �*�=��\$�D$d�L$�D$h�L$�\$ �D$l�L$�\$$�U�E����M�U�D$ ���\�E�M�D$$���\�U�E���D    ��O�QH��$0  SP�RH��   ��$�   �ل$�   ،$�   ل$�   ،$�   ��ل$�   ،$�   �������������@t���D$0    ����D$,    �3�=��\$ل$�   �L$ل$�   �L$�\$,ل$�   �L$�\$0�M�U����E�M�D$,���\�U�E�D$0���\�M�U���D    ��O�HH��$�  SR�QH��   �|$x�ل$�   ،$�   ل$�   ،$�   ��ل$�   ،$�   �������������@t���D$<    ����D$8    �0�=��\$�D$|�L$ل$�   �L$�\$8ل$�   �L$�\$<�E�M����U�E�D$8���\�M�U�D$<���\�E�M���D    �D$��t-�U�E �M���U�E$�M���U(�E��D$��t�E�ES�������؅�����_^][�İ  Ð��������������D$�T$��8  SUV��$H  3ۉF��$T  W��^�^�^�^�V�F �^�]�  ;�t�F��O���   ���R(;�u�FhD���h�   P�k�  ��;ÉF�  �NS��QP���  �VhD���h�   R�9�  ��;ÉF��  �NS��QP��  �VhD���h�   R��  ��;ÉF��  �F�NS��PQ��  �F��hD��@h�   R���  ��;ÉF�o  ��z�  ��;��k  3�O���   ���R=G  ��  �FhD�h�   jD�<(�|�  ��;�t�N �VQ�NR�VQ�RWQ���:����؅ۋV�*��  �F�L$Q�ˉ(舊������   h����$�   ��  ��O���   ���PxP��$�   Q��$�   R舷  P��  ����$�   ��  ��$�   �׶  h����$�   薶  ��$�   P�y�  ����$�   誶  �L$Q�L$L�l�  �T$HR�R�  ���L$H�  j ���-�������  h����$�   �4�  ��O���   ���RxP��$�   P��$  Q�ζ  P���  ����$  �)�  ��$�   ��  hl��L$l�ߵ  �T$hR���  ���L$h�t  ��O���   ���R=�q �^  �F�<(��O�Q@SW�Rt�؃�����  W���z������  ��O�H@W�QhP�T$R�p��������   h����$�   �J�  ��O���   ���RxP��$�   P��$0  Q��  P��  ����$(  �?�  ��$�   �3�  hL���$�   ��  ��$�   R���  ����$�   �  ����~���؅�u|h����$�   踴  ��O���   ���RxP��$�   P��$   Q�R�  P�|�  ����$�   譴  ��$�   衴  h,��L$�c�  �T$R�I�  ���L$��   �D$P���!�����uqh���L$,�/�  ��O���   ���RxP�D$,P��$   Q�˴  P���  ����$  �&�  �L$(��  h ��L$<�߳  �T$8R���  ���L$8�w�F�(�th���L$\足  ��O���   ���RxP�D$\P��$@  Q�R�  P�|�  ����$8  譳  �L$X褳  h���L$|�f�  �T$xR�L�  ���L$x耳  ��O���   ���R(��3ۃ�;������_��^][��8  � h���XH����_��^][��8  � ������SV��F3�;�t	P�M�  ��9^W�^t'�F3�;�~�F��;�t�j��F���FG;�|�F;�_t	P��  ���F;É^t	P���  ���F;É^t	P���  ���^^[Ð������������VW�|$��t�q3���~�Q9:t@��;�|�_^2�� �I�����T$�t���@R  ��t
_^�   � _^3�� �����������V��FW3���~!�F����t�F���P�P�R�FG;�|�_^Ð��������������VW���G3���~�G����t��R�GF;�|�_^Ð��������S�\$�U�l$�h�V�t$W�z�   ��K�H��C�B��A��O�JHj h�  P�Qx����tE�����  ����t8��O���   ���P=�q t��O���   ���R=G  u��p�s��A��O�JHj h  P�Qx����t��B�C����  ��t�C��tU��u�{tJ�D$ ��uB��O���   ���R=�  u+��A��uh�Ih���|  _^]�   [� Q�Q��_^]�   [� ��������������D$��(V��L$4hD�h�  j0��N(�l�  3Ƀ�;���   �H�H��H�H�H�H �H�H�H,�H(�H$W���Љ:�z�z�L$�D$  �?�T$�P�щP�P�L$�P�L$�D$  �?�T$�P�щL$�P$�L$�L$�P(�P �D$  �?�T$�L$�L$�L$�P,_�3�Q�T$ Rj�F�D$Dh   @�F�Q�L$4�L$8�L$<P�L$(�D$(���t$4臮  ��^��(� ��������������hD�hF  j�_�  ��Ð�����������D$��tP�r�  Y� ���������������D$��L$��P�Q�P�Q�@�A� ���������������V��F��t	P� �  ���F    ^Ð�����O�I���   �Rx�L$jh�   Q��謰  �� ���������OSUVW��~�HHj h�  W�Q|�\$ ��F��O�BHh�  W���   �L$,��F��O�BHj h�  W�P|�l$<�E �F ��O�QHh�  W���   �L$H��F$���(��t �}  t�D$�8 t�9 t_^]�   [� _^]3�[� ������������������  SUVW�ًC��O�QH3�Wh'  P�Rx��;ǉD$<u_^]2�[���  � �s$�v��P�s�  ��;�tN;�|�H�V�y�9�y���Ju�D$D��|$D9{$�|$�?  �L$D3�L$ �s �L.�D.�{�;��uz�@�D����I�d���Q�$Q�@�a�$Q� �!��$�   �$��
  ��v�@��$�   Q��P�v��R��$�  P��  ��P��$8  Q��
  P��$�   R�Z�I��R�@��Q��$,  R�  ��P�F�v�@��Q�v��P��$H  Q�r  ��P��$P  R�
  P��$�   P�
  �L$4��$�   �щ��$�   �B��$�   �B�D$0����@�L$ �K$��;��D$�����3��C$����$�  �O  3��O��$�   PǄ$�       Ǆ$�       Ǆ$�       Ǆ$�       Ǆ$�       Ǆ$�       Ǆ$�       Ǆ$�       Ǆ$�       Ǆ$�       Ǆ$�       Ǆ$�       �QD�L$@WQ�R<ل$�   �C �(ōI����ل$�   A����ل$�   �\��Hل$�   �I��Aل$�   ��ل$�   �\��Hل$�   �I��Aل$�   ��ل$�   �\��@ل$�   �@��@ل$�   G��ل$�   �\��C$;��������$�   �p�  �S$�C �Kj RPQ��$�   ��  ��u��$�   �v�  _^]2�[���  � �C3Ʌ��L$ �.  ��$�  +Ɖ�$�   ��$�  +Ɖ�$�   ��$�  ��+ƉL$�l$@�D$<��O3��D$l��$�   �Bx��$�   R�T$pRQ��$�   Q�P�����$�   ����������~/�L$l�׋�l$D�@�D� �D� �Ƀ�J�@�����@��uۋl$@�������������������������@t"���D$,    ���D$(    ���D$$    ���"�=��T$���\$$���L$�\$(�L$�\$,��$�   ����D$$�T$H�T$,�����T$������L$(�T$����E �M�T$�U�l$@�D$`�D$�T$h�S�L$d����$  �A�I��$  �E ��$  �M�D$8    �D$4    �D$0    �D$P    �D$L    ��$�   ��$  ��  �D$l�D$0�D$��$�   �L$�	�C ���|ȋA;�����������Q  �D$|�;D$ �/  �@���<�/��$�   ل$�   ؤ$  �o���$   ل$   ؤ$  ��$  �l$@ٜ$�   ل$  ؤ$  ٜ$�   �0ؤ$�   �\$�D0ؤ$  �\$���L$ل$�   �L$ٜ$d  ل$�   �L$ٜ$h  ���D$4؄$d  �\$4�D$8؄$h  �\$8�L$ل$�   �L$ٜ$p  ل$�   �L$ٜ$t  ���D$L؄$p  �\$L�D$P؄$t  �\$P�D$�L$���D$�L$���D$�L$�D$|��H�D$|������L$��$�   ��H�L$��$�   �f������T$���T$H���\$0�\$�\$�Ɋ�$�  ����  ���������D$L�L$ٜ$�  �D$P�L$ٜ$�  �D$0�L$�D$4�L$ٜ$�  �D$8�L$ٜ$�  ��ل$�  ؤ$�  ٜ$�   ل$�  ؤ$�  ٜ$�   ���L$$ل$�   �L$(��ل$�   �L$,�����L$$�\$p�D$(���\$t�D$,���\$x���d$pل$�   �d$tٜ$X  ل$�   �d$x����ل$X  ،$X  �����������������@t)���D$\    ���D$X    ���D$T    �,����������=������\$Tل$X  ���\$X���\$\���D$X��$�   �L$$�T$T�D$(�D$X�L$T͉�A��T$\Q�Q�$Q�D$4�L$\�D$d�L$,���$Q�D$h��$�  �L$4�D$d�L$8���$��  �D$<��$x  ��$|  ŉ��$�  �P�H�v  �D$PQ���$Q�D$T���$Q�ɍ�$H  ���$���  �D$8Q�L$�$Q�D$<�L$�$Q�D$<��$T  �L$�$�j  ل$P  Qؤ$H  �$Qل$T  ؤ$H  �$Qل$T  ��$�   ؤ$H  �$�(  �D$8Q�L$�$Q�D$<�L$�$Q�D$<��$<  �L$ �$��  �D$PQ�L$�$Q�D$T�L$ �$Q�D$T��$0  �L$$�$��  ل$,  Qؤ$<  �$Qل$0  ؤ$<  �$ل$,  ؤ$8  Q��$$  �$�  ل$�   �L$`Qل$�   �L$l��ل$�   �L$h���D$l���$Q�D$l���$Q��$�   �L$l�$�9  ل$�   Qؤ$�   �$Qل$�   ؤ$�   �$Qل$�   ��$�  ؤ$�   �$��   ��$�  R��$�  P�B  ل$   �L$h�ل$(  ��$�   �L$p͉�P���Qل$$  �@�L$l���A�L$`��QQ��$�  �$R�[  P��$(  P��$�  Q�u  P��$�  R��   ��L$\�� ͉�P�Q�@�A�L$ �|$�CA����;ȉL$ �|$�l$@�	����L$DQ�n�  ����$�   ��  _^]�[���  � �T$���L$��L$�P�H� ��������L$�D$��H�A����A��@�	���A�H�A�H�D$����X�XÐ�����L$�A�A��������������������������������@t�D$��3ɉH�H���=��D$�T$�I�D$�I�D$�	��X�XÐ�������D$�D$�H�D$�H�D$��D$��X�XÐ�����������D$�@�L$�a�@�a� �D$�!��X�XÐ������������0��V�p�D$8W�   �|$��D$��T$�L$�P�T$ �P�T$$�P�T$(�P�T$,�H3ɉP �T$0�H�H�P$�T$4�H,�L$�P(�T$�H0�L$_�P4�H8�@<  �?�^��0� ���������D$�Q�I(PR����� ��������������0  �D$0P�P�����u�D$0�L$0Q�L$��  Ph���L$�۟  P�T$(R萠  P躰  ���L$ ��  �L$ ��  �L$�ܟ  ��$8  P�L$$蛟  ��$4  PQ�L$艟  P�T$R�>�  P�h�  ���L$蜟  �L$ 蓟  �L$ 芟  ��0  � ���xU��E��O�Q@P�Rh�M ��$�   ��h#  Q�� N  R����  ��u	2�]��x� ��O�QHS��$�   ��VWPt1�D$,P�RH��   �|$0�L$0�T$4�D$8���L$�T$�   �D$,P�RH��   �|$0��D$T�L$T�D$X�L$X���D$\�L$\�������������@t���D$$    �D$     �D$    �&�=��D$L���\$�D$P���\$ �D$T���\$$�؋L$�T$ �D$$�L$�T$�D$��$�   ����   �ۋu�   �|$(�t�D$0    �D$,    �D$(    �L$(Q�T$\R��T���D$ �H$���D$�H���D$�H��� �\$�D$�H(�D$�H���D$�H���@�\$ �D$�L$ �H,�D$�L$�H ���D$�H���@�D$�D$�\$$�T$$�T$��$�   �D$�L$��T$_^[�H�P�@  �?�]��x� ��������SV��F��u^�[��ÍL$�A�  j �D$P�L$ Q�L$�D$$�  �D$(    �D$,    �4�  �NP�+�  ����ۍL$���J�  ��t"h�Ih���������L$�<�  ^�[��ÍL$�;�  ���L$����  ^��[��Ð������0h'  賸  ��P�L$�6�  �L$ ��  ��u�L$ 耜  �   ��0�Vh$��L$(�8�  h��L$�*�  j �D$(P�L$Qh�� j�T$RhIr �ؼ  ���L$���*�  �L$$�!�  �L$��  ��^��0ÐVh0�jj��  ������t����  �����^�3�^Ð��VW�|$��j ��蟰  � -�  tUHt!�D$�L$�T$P�D$QRWP���Ƿ  _^� ��O�D$�Q@P�Rh����tj h�  ����  ��u_3�^� _�   ^� ���������O�����4!  }*h���L$��  �L$ Q�v�  ���L$ �*�  3�����O  �j�����u����,  ��u�����d����u�����W������؃�Ð����������X���F.  �������D$�� tHt3�ù�O藵  �����ø   Ð����������D$SV�t$W�   �κ   ������Ju��Ou�_^[Ð��D$�L$$�D$�L$ ���L$�D$�L$$�D$�L$ ���L$���D$�L$�D$�L$���L$��Ð��������V�t$�F<�N8�V4WP�F,Q�N(R�V$P�FQ�NR�VPQR�����|$4��F<�N8�V4P�F,Q�N(R�V$P�FQ�NR�VPQR�R������_�F<�N8�V4��HP�FQ�NR�VP�FQ�NR�VPQR�!����_�F,�N(�V$P�FQ�NR�VP�FQ�NRP�VQR��������_�F<�N8�V0��HP�F,Q�N(R�V P�FQ�NR�VPQR��������_�F<�N8�V0P�F,Q�N(R�V P�FQ�NR�PQR�����_�F<�N8�V0��HP�FQ�NR�VP�FQ�NR�PQR�i������_�F,�N(�V P�FQ�NR�VPQ�F�NR�PQR�<����_�F<�N4�V0��HP�F,Q�N$R�V P�FQ�NR�VPQR�����_ �F<�N4�V0P�F,Q�N$R�V P�FQ�NR�PQR��������_$�F<�N4�V0��HP�FQ�NR�VP�FQ�NR�PQR�����_(�F,�N$�V P�FQ�NRP�V�FQ�NR�PQR�������_,�F8�N4�V0��HP�F(Q�N$R�V P�FQ�NR�VPQR�V������_0�F8�N4�V0P�F(Q�N$R�V P�FQ�NR�PQR�)����_4�F8�N4�V0��HP�FQ�NR�VP�FQ�NR�PQR��������_8�F(�N$�V PQ�F�NR�VP�FQ�NR�PQR������W<�F��H�O�����G�N0���F �O���=���������O�_���O�_���O�_���O�_���O�_���O�_���O�_���O �_ ���O$�_$���O(�_(���O,�_,���O0�_0���O4�_4���O8�_8�����_<_^��Ð����D$�L$� �	�T$�@ �I���@�I���A�H0����@�I�@$�I����H���@4�I���Z�@(�I�@�	���@8�I���@�I���Z�A�H<�@�I���@,�I���@�	���Z�@�I�A����A�H0���@ �I���Z�@�I�A�H���@4�I���@$�I���Z�A�H�@8�I���@(�I���A�H���Z�A�H�A�H<���A�H,���A�H���Z�@�I$�A ����A,�H0���@ �I(���Z �@�I$�A �H���@4�I,���@$�I(���Z$�A$�H�@8�I,���@(�I(���A �H���Z(�A �H�A,�H<���A(�H,���A$�H���Z,�@�I4�A0����A<�H0���@ �I8���Z0�@�I4�A0�H���@4�I<���@$�I8���Z4�A4�H�@8�I<���@(�I8���A0�H���Z8�A0�H�A<�H<���A8�H,���A4�H���Z<Ð�����������Q�T$��3ɉ�H�H�H	�H
�H�P�H�H�HYÐ�������SVW���_�w;�t�j �����(;�u�OQ�I�  ���G    �G    �G    _^[Ð���������������   SUV��W�\$4�  ��$  ��u���h��P��  �������|$uj��$  腩��_^]2�[���   � W�   U�D$8jP��  U�L$Dh��Q���  ����Wt>�@�  ��$  �����t  �A����_  <��W  _^��]�A�2�[���   � j��$�   j|R��  ��$   ����t�C	�    ��$�   t��v�C
��$�   ���   ��$�   =DXT1tk=DXT3tU=DXT5t?W��  ��$  ������  �A�����  <���  _^��]�A�2�[���   � ��  �k�C�~��  �k�C�o��  �C   �C�\��Au��$�    u���  �C �k�>��@�i�����$�   �� u��  �C �k����E������  �C �C   ����$�   ��$�   ��l$(�|$<�t$ �D$    �t$ �K���D$`� u�D$�� �K	���D$$    Ƀ�A���`  ���D$8�����D$@�����D$,��t$ �l$(�|$<WU���T$$��PVWU�L$l��  �T$�D$lRPj�L$h�  P���  ���L$\Q����  �C	��u0��$  ��t%�T$l�D$h�L$dR�T$dPQR�L$l�Y  P����	  �l$8���   �t$@���   �|$,���   ��$�   ���D$tH�D$�D$���D$    ��   ��u����   VU���T$$��PWVU�L$T�  �D$�L$TPQj�L$P��  P��  �C	����u0��$  ��t%�T$T�D$P�L$LR�T$LPQR�L$T�  P����  �L$|�D$DPjQ��$�   �q  �����   �����   �����   �L$D�7  �D$�L$@;��D$�0����K�S�s+Ѹgfff��������Ѓ�����   �F��t+ȸgfff��������у���w�   ���.  ��݋�y3�����R�H�  ����FUWP���6  �L$\QjP�ΉD$�c  �T$�F��(RPW���  �N�VQR���P  �FP�W�  ���T� ���ΉV�  �\$4@���L� �N�n�   ��+׸gfff��������Ѓ�sN�W(RQW���  �n�D$\P��+ϸgfff��������Ѹ   +�PU���  �V�L$\QRW�I  ���-QQ���Q���W  �FP���PW�Y  �D$hP�O(QW�  ���F(�L$\��  �D$$�S	@�ډD$$҃�B;�������D$P��  ��$  �����Ct)�A���t<�t_^��]�A��[���   � IQ�,�  ��_^]�[���   � IQ��  ��_^]2�[���   � �SUV���F    �    �F �F	 �F
 �F �^�nW��;�tW����  ��(��(;�u�^;��t�j �����(;�u�_�n^][Ð��������������SUV��F��W��   ��I��uh���������Iu_^]2�[Ë~���q  �O�P�GPj QRj h�  ��I3�3ۋ~�G����   �O +ȸ���*���������;���   ��;E�  �L;�T;P�Qj RPUh�  ��I��맋~�����  �OPh  Sj QSj h�  ���3�3�N�A��tK�Q +и���*���������;�s1�y�/C�  ��T/P�Fh  Qj RPSh�  ������_^]�[Ð�SUV��F��W��   ��I��uh��������Iu	_^]2�[� �|$�^�<�����|$�   �L�TP�DP�j Q�L$(RPj Q��I3�3ۋV�D�����   �Q +и���*���������;���   �y�;E�  �L;�T;P�D;Q�j R�T$(PQUR��I�|$��뚋|$�^�<�����|$�{  �L�TP�h  P�Fj Q�L$,RPj Q���3�3ۋV�D���tT�Q +и���*���������;�s:�y�;E�  ��T;P�D;h  Q�Nj R�T$,PQUR����|$���_^]�[� ������h��  j �d�������Ð�������������VW��3����  PV���;�����tF��|�_�^�_2�^Ð������QSU�يC��VW��   ��I��uh4��������Iu_^]2�[YËs���O  �N�VP�FP�Fj Q�RPQj ho�  ��I3�3��k�E���  �U +и���*���������;���   �uA�L$�7��  �L7�UP�D7Q�L7�t$j R�PQRVho�  ��I�΃�딡�I��uh$��������Iu_^]2�[YËs���  �N�VP�h  P�Fj Q�KRPQj ho�  ��I3�3��s�F��tU�N +ȸ���*���������;�s;�v�7E�1  ��T7P�D7h  Q�L7j R�SPQRUho�  ��I���_^]�[YÐ�����������D$�L$S3ہ��  �Ã�������K������؍A��������[� ��A�D$�D$� �A��<��SV��   �A
����   �A	����   �\$H�A�S�s��   ����������L$9C��   �KPQVR�L$,�{  ���4  �L$�D$�'  �s���D$�D$    ~fUW�T$�C�T$P����K�l$���3҅ɉD$ ~0�t$P�������ȋD$���|$P�K�D$ �B;щ|$P|ЋD$�s@;ƉD$|�_]�L$Q���  �L$�
  ^[��<� �SU��E��VW��   �D$$�t$ ����\$�ș�����L$ ���  �Ë\$���D$�\$�t$$��+���~)�D$WSV���  �D$�+�H�D$u�L$ �D$�\$�T$$�J�\$�T$$u�_^][� �D$���ȋD$���U �������  �L$$t(JtJ��   �   �D$�� ��   �D$�� ��   �D$�� ��������~Q�|$���މt$ �p������T$��L$$QW���T$$�D$$PV���T$$SWV���%   �L$ �D$��H�D$u�_^][� �����������S�\$UVWS袜  �T$�ˋ�������͋l$�����ˋ������ʃ����������ʃ�P�躜  ��_^][� S�\$��W��~.�D$V�pj�NQV���~���j�VR�FP���m�����Ku�^_[� ����D$��SU�l$�ىl$��   V�M�UW�}�u�L$ �T$���D$�D$jWP������jVU�������T$�D$�   ���T$�T$ j��P��V�ˉD$�T$,������L$ jWQ��������T$�L$ �   ЉT$�T$������D$H�T$�L$ �D$�k���_^][��� �����������V�t$ �N��f��@�D$    f�T$���D$�D$�T$���Ѐ��T$	�D$���Ѐ��T$
�D$���Ѐ��D$�T$���Ѐ��D$�T$���Ѐ��D$���T$�D$������$�T$�D$����f��@�D$    f�T$���D$�D$�T$���Ѐ��D$�T$���Ѐ��D$�T$���Ѐ��D$���T$�Ѐ��D$���T$�Ѐ��D$�T$���ЉD$��$�D$���T$�D$�T$%�   �����   T$�����   T$�����   T$�����   T$�����   T$�����   ����   �T$���   �D$�L$
�T$	%�   �����   ��L$�����   T$�����   ��L$�����   T$�����   �������   T$����   �����   ^��� �����Q�D$��V�t$�L$�t$~wSUW�n�^�~���D$�D$�L$P�����L$j����V�L$ �L$��W����������L$jSU������T$�D$����������H�T$�D$u�_][^Y� ��������������V����  �D$t	V諘  ����^� ���D$�T$VP�D$��L$QRP���b  �L$3��F�F �F$�N����^� ������SU�l$$VW��U�|$(�i  �D$,3ɍw��N�N�N���L$�L$�E;��  �M +ȸ���*��D$�������;���  �L$�]�VًN+Ѹ���*��������Ѓ�����   �n��t��+ո���*��������Ѓ��T$w�D$   ��u3��+͸���*��������ыD$��D$}3��@��Q�	�  �D$$��F��;ǉD$t"��D$PU�8  �D$������;ǉD$u�SjU���h	  �V��URW���	  �F�NPQ����  �VR� �  �D$ �|$$�@�ǉN�����u  �l$,@�@�׉F�~�   ��+׸���*��������Ѓ�sS�WRQW���  �n��+ϸ���*���������S�   +�QU���  �VSRW�	  �F�l$8�����F�2QQ���Q���U  �FP���PW�	  S�GPW�L	  �F�����F�L$�D$�|$$A���L$�D$3��������_^][��� ��������D$SUV��;�W�t$�  P�  �n �^����;�tW���j  ����;�u�n;݋�t�j �����;�u�3��^�D$�|$(�D$�G����  �O +ȸ���*��D$�������;���  �_�D$�N�V�+Ѹ���*��������Ѓ�����   �F��t+ȸ���*��������у���w�   ���  ŉD$ y3��@��R蚔  ����FUWP����  SjP�ΉD$(�  �L$�V��QRW����  �F�NPQ���v  �VR譔  �D$$�@�L� �N�����%  @�@�D� �F�n�   ��+׸���*��������Ѓ�sF�WRQW���[  �n��+ϸ���*���������S�   +�QU���r  �VSRW�7  ���)QQ���Q���  �FP���PW�G  S�GPW�  ���F�L$�D$A�L$���A���_��^][��� �D$_^][��� ������SUVW�����o �_��;�tV���@  ����;�u�o ;݋�t�j �����;�u�_ �w;�t�j �����;�u�GP�\�  3����ωG�G �G$�W  _^][Ð�V���H  �D$t	V�+�  ����^� ���D$�T$V��L$P�D$QRP�����F    �%  ��^� ���������������3�S��V�t$�C�C�C�C�C��9FtF�F�C�N�K�V�K�S�FWQ�C�:�  �C�N�v���������ʃ��_^��[� ^��[� ���������������SV�t$��;�tR�   �F��tF�F�C�N�K�V�K�S�FWQ�C�Ƒ  �K�щC�v�������ʃ��_^��[� ^��[� ��������������U   ������AÐ�����������V���8   �D$�L$�T$�F�D$P�N�V�F�F�  ���F^� ������������V��FP脑  ���F    ^Ð��������A��uËI+ȸ���*��������Ћ�Ð��������������V�t$W�|$;�t�j �����;�u�_^� ��������������V�t$W�|$;�t�j �����(;�u�_^� ����������������SU��MV�u+θ���*��������W�|$ �;׉l$�s  �]��t��+˸���*���������;���r�υ�u3��+󸫪�*��������Ѝ
���D$ }3��@��Q���  �u�T$ ��;�D$��t��tV���V����T$����;�u����v���t�T$$R���0�����Mu�T$�t$�N���;э,�L$t&��+�+���tV��������L$����;�u�t$�^�v;�t�j �����;�u�L$�QR袏  �D$$�t$�L$�@�ƋA�����Qu3���_�։q^]�A[��� �Q+и���*�����������_�։q^]�A[��� �\$��+˸���*���������;���   ���;ލ�D$�L$ t$��+��t
U�����L$ ����;�L$ u�l$�u��+˸���*���������+�t��t�L$$Q���������Ou�};ߋ���   �T$$R���6�����;�u��q��vt�����+�;���D$t��tW�������D$����;�u�l$�}��+�;�t����V�������;�u�D$�4;�t�|$$W���������;�u�D$E_^][��� �����������S�\$V�t$;�t#W�|$��tV����������;�u��_^[� �D$^[� �������D$��v"S�\$V�t$W����tS��������Ou�_^[� ����A��uËI+ȸgfff��������Ћ�Ð��������������S�\$V�t$;�t#W�|$��tV���������(��(;�u��_^[� �D$^[� �������D$��v"S�\$V�t$W����tS��������(Ou�_^[� ���V�t$W�|$;�tS�\$S���u�����;�u�[_^Ð���������S�\$V�t$;�tW�|$����V���?���;�u��_^[ËD$^[Ð�������������V�t$W�|$;�tS�\$S���e�����(;�u�[_^Ð���������S�\$V�t$;�tW�|$��(��(V���/���;�u��_^[ËD$^[Ð��������������L$��t
�D$P����Ð�������������TX���u
ȈTX�   �������h@� �/�  YÐ����� V�t$(W�D$3�P�Ή|$������uh�Ih����� ���_^�� �SU�L$,Q�T$$R�D$ P�L$(Q�Ή|$,�|$03�|$$�|$8�{�����uh�Ih������  �5��ht�  �֋T$RWh  j����D$�@��P越  ���D$�@��Q褊  ��D$ �@��R蒊  �D$ �D$$�@��P�~�  �����؉\$(�q  ���i  �D$���]  ���U  �L$��R�L$4P�D$SPUW�v�����uh�Ih���1  hu�  ��Wj h  ���h��  �dJhx�  ��S���j h  j��h��  �dJhx�  ��Uj h  j��h  �dJhx�  �֋L$Qj h  j�ӋL$�qE�����j �D$(P���Rx��}h�Ih���   �L$�D$4�P�R��tG�D$$3ۅ�v3�S���R|��|<�D$ �L$,Ph  ��    Rj����D$$C;�r͋�����   �L$��R�1�L$4h�Ihl�������L$��R�h�IhP��L$<������5��ht�  ��hu�  ��h  �dJhx�  ��h��  �dJhx�  ��h��  �dJhx�  �֋D$(P���  �L$Q��  U��  W�߈  ��][_^�� Ð���U������0VWh  �?j j j �l�h A  �đ�5ȑh  �֋=̑��h   ����h  �?j j j j j j j �p�j�t��5x�h  �j h  �j ��h  �j h  �?j ��h  �?j h  �?j ��h  �?j h  �j ���|��E�Mhp
PQ�L$�H����L$�����_^��]Ð��������V���8�  �D$�F�F%'  ����^� ������������������IVj ��P�L$Q���D$&'  �D$    �x  ��Ij R�D$P���D$('  �D$    �ax  ^��� �����������D$��D-&'  V����   Ht4H��   ��IP�L$�D$('  �D$    Q���y  ��us^��D� �L$,�+g  j j j �L$8�g  ��tG�T$R�L$0��g  ��IP��o  �L$�o  ��Ij P�L$Q���D$&'  �D$    �w  �L$,�Hg  �   ^��D� ��IR�D$�D$&'  �D$    P�U��������������Vh �jFj���/�  ����t
V���`���^�3�^Ð����������L$��t�j�� �����������������xVh �jSj�.n  ����t���Pn  ����Iu^��x���I    3�^��x�h �jWj��m  ����t;���n  ����Iu7��I��t���{n  V��m  ����I    3�^��x���I    ��h �j^j$�G�  ������t���7�  �$����3ɉ�I������Iu^��x�h'  ��  ��P�L$�m  �L$�sn  ��u�L$��m  3�^��x�j j �L$Q��Ih�q ��  ��u�L$�m  3�^��x�h���L$�tm  �T$R�L$d�e  P�D$HP�i  ��P�L$0Q�}f  ���L$D�Ae  �L$`�8e  �L$�_m  ��f  ���D$tGh1D4ChCD4Cjjj�T$<R���g  ��t'��I�L$P�g  ��t��IQ�L$�g  ��uNh�I�L$��l  ��I�T$R�m  �L$��l  h|��L$�l  ��I�D$P��l  �L$�l  �L$Q�cf  ���L$(�wd  �L$�l  �   ^��xÐ�����hh���L$�Ol  �D$P�L$P��c  P�L$4Q�h  ��P�T$R�Xe  ���L$0�d  �L$L�d  �L$�:l  ��e  ���D$ tPh1D4ChCD4Cjjj�L$(Q����e  ��t#��I�L$ R�}g  ��t��I�L$ P�jg  �L$ Q�e  ����I��t��I�P�R��I��t	P��  ����I��V��I    t���k  V��j  ����I����I    t���vk  V��j  ���L$��I    �*c  ^��hÐ�����D$��Ijh�   P�)m  �Ð�������I��   VP�L$ �j  h���L$��j  j �L$Q�T$R�L$(��k  �L$����j  �D$P�L$@�~j  ����   h���L$�j  ���Ak  �L$���j  �L$�-k  �ȋD$+�+�Q�V�T$4R�L$(��k  P��$�   P�L$dQ��l  �T$$��PRj �D$|P�L$0�k  P��$�   Q��j  ��P�T$R��j  ��P�L$@�lj  �L$�3j  �L$|�*j  �L$l�!j  �L$\�j  �L$,�j  h���L$��i  j �D$P�L$Q�L$H��j  �L$����i  �T$<R�L$P�si  ����   h���L$0�i  ���6j  �L$,���i  ��$�   P�L$�ji  �L$<�j  �ȋD$+�+�Q�V��$�   R�L$H�j  �L$P�D$PQj �T$|R�L$P�j  P�D$hP��i  ��P�L$4Q��i  ��P�L$P�ai  �L$,�(i  �L$\�i  �L$l�i  �L$|�i  �L$�i  h���L$��h  �T$LR�D$P�L$4Q�ri  ��P�L$ �i  �L$,��h  �L$��h  ��$�   jh�   R�L$(�j  �L$L�h  �L$<�h  �L$�h  �^�Ĉ   Ð������Aj?j P��r  �����Ð�����������V��NW��  ����u_�   ^ËW���P(�W���R,����r  _^Ð������������ �������������3�V���F�F�F� ��F��^Ð���D$�T$SV��L$3ۉN�NH��^�F�V<�F@����^D�����^P�^T�^X��^[� ����������������SUV��nHW���m����~L3�;�t�������W�~  ���FDP�^L�~  �~T��;��^Dt���$���W�~~  ���~X;��^Tt���Z4��W�d~  ���~P;��^Xt������W�J~  ���;É^Pt@9Xt;�@;�t(SP�ԑ��A;�tP�ؑ��P�@RP�PO��QR�TO� ��+A�D$�\$�l$���T$ �@��$h��R躙  �D$(P������������_^][��Á�   SVWj���>}  ����t	���P����3����u
h���  ��$�   ��V<R�����F�F<P�������F�@�L$�D$�~�P��H��j�  ���F@��P��|  �����FDu
h���J  �V<UR�����F�F<P�����N<Q�F������V<R�F �����F�n ���F�ŉD$ �~$�D$ �����  +��~�|$ �؉^,�D$ �^8���܌  �؉F0ÉF4�F<P�)�������]u
hh��  �N<Q�N�������u
h@��  j�|  3���;�t�V�NRQ�������3�;ǉFLu
h��l  �V<PR�NH������u
h ��Q  �N�   �D$8�D$H������   %A   �D$L����D$P�L$Q��T$`S�T$(R�D$4�D$,    �D$0    �D$4-   �\$8�D$<   �D$@'   �D$D   �D$L   �D$P   �D$T"   �\$`�D$dB   �|$l�PR�dO;���  9|$��  �N�V�D$P�D$Q�R�|$�PR�HO��A��B;�u
h���^  P�LO��A��B;�u
h���?  P�X���A��H;�u
h���   �PQR�ԑ��u
h`��  �F�NPQWW���h  �?WWW�l�9~t�  ��th  h4�  �h�WhX��S  ����}
h0��   j0�z  ��;�t�V<R��胣���3�;ǉFPu
h��   j,��y  ��;�t�N�VPQ�R�R���\-���3�;ǉFXuh���Mj$�y  ��;�t�NX�VQ�NPR�V<QR�������3�;ǉFTuh���_�^^��[�Đ   � h��������_^2�[�Đ   � ���������V��F��u3�^����F�F���`�����Au�`������\$�����`��D$�X�����Au�X��������X�� ��q�  � �P�e�  �NLP�|���^��Ð��������V��F��Wu_�   ^��ËF0���D$t6�V,�N8�F +ʋV$+��ʉL$�D$�F<�D$���t$�D$�v�$P��F$�N<���v�$Q�����VT�F<�NX��RP�1����H�PQR�ԑ��u
h��   �NT�����FX�NT�V<PQR����������NT�&����FD�N�VPh  h  QRj j �d��F3���~�VD�NL���F@�PW�H����FG;�|�NLQ�NH������uh���������F �V8�NB�ɉV8��u_�   ^��Ë~43�;���_^J����Ð��������������T$���P�T$�P�T$2ɉP�T$�H�P�H� h�� �V���   �D$t	V�kw  ����^� ���h�Ð���������AÐ�����������V��F���FtW�=Аjd�׊F��u�_^Ð�������������D$�T$VP�D$��L$QRP���B����p���^� ������V���   �D$t	V��v  ����^� ���p��U��������QV�D$Pj ��Vh�j j �D$    �F�Đ��uhD��F�8�����2�^Y�P�Ȑ�^YÐ���UW�)  ��uh�������|$�O���\  ��   �b�  j Pj j h�   h�   j j h  � h��h��j�����uh�������|$�O���  �}Vj\�}u  �|$����t�O�WQ�ORQ����������uh���o����O����  �2SU�����uEhh��L������O�  ������V�tu  ��[U���^�OQ�������G _3�]� P��������t��G3ۄ�u���u��������؃�t��V0�N,�F8j B+�RP���c����OP��  �G��t�뀐�D$�T$VP�D$��L$QRP���2����L$�N�x���^� ���������������V���   �D$t	V�t  ����^� ���x��5��������QV�D$Pj ��Vh�!j j �D$    �F�Đ��uhD��F������2�^Y�P�Ȑ�^YÐ������   SV�c�  3ۋ��\$,�\$ �\$� ��D$<��  ��uh����������i  SVSSh�   h�   SSh  � h��h��j��;ÉD$0uh���������(  UWP���;ÉD$u
hh��S  ��$�   �M��  �M���t$ ��  ���EP�|$�����M��Q�\$ ��������ۉD$u��u��u���  �D$3�3��t$�D$�D$ ������������Au������� ��H�  ���؋������� ��1�  ���؋�+�v�L$�D$�D- +��P��H���  ���D$<��P�dr  �����D$u
h���`  j�Hr  ����tWV���h������D$ uh��7  �D$     h��%  ��$�   �K���ڽ   �   �D$\�D$lҁ�A   �����T$p�L$Q�T$DR�T$U��$�   �D$8P�L$XQR�D$D    �D$H    �D$`-   �l$d�D$h   �D$l'   �D$p   �D$x   �D$|   Ǆ$�   "   ��$�   Ǆ$�   B   Ǆ$�       �dO;��U  �D$���I  �L$@�T$�D$PWVQR�D$(    �HO���D$4u
h���  P�LO���l$(u
h���  U�X����D$$u
h����  PU�ԑ��u
h`���  WVj j ���h  �?j j j �l��C��t��  ��th  h4�  �h�j hX���I  ����}
h0��y  j0�ap  ����t�KQ���ϙ�����D$uh��N  �D$    h��<  j,�$p  ����t'�S�L$R�T$QR���#�����D$uh���  �D$    h����   j$��o  ����t+�L$�SQ�L$R�SQR���������D$uh���   �D$    h���   �L$P�CP��(���L$$QU�ԑ��u
h��   �l$���V����T$�CRUP�������������w����l$Uh  h  WVj j �d�3���~�L$ UV�����L$<F�;�|�KQ�L$$j�j*�����KP�F  �h���
������t$ 3�;�t���V���V�0o  ���T$R�#o  �t$��;�t��豤��V�o  ���t$;�t����$��V��n  ���t$;�t��聙��V��n  ���|$4;�t.�t$(;�tSV�ԑ�D$$;�tP�ؑVW�POW�TO�D$8P���_]��$�   �NQ�������� �+D$<�D$$�\$(�l$$����$�   �@��$h��R�<�  ��$�   P�!������F ^3�[���   � �������������V����a  �   �F�F3��F�F ����F(�F,�����F0����*}  �F��^Ð��V���   �D$t	V��m  ����^� ��V��F��W�~���t+��O�QPj P�RL����t�FP�F  ��W��|  �����ja  _^Ð��������   V���c  h�  ���Vb  �F�NPQj j ����a  �~(�u3h�  ���1b  hp��L$��U  jj�T$R���3b  �L$��U  �F���1  ��O�QPP�RH�����  �F��W��   ��O�QP�R��O�Q���FP�|$�R�����D$��   ����   �F���D$��   �F���D$��   �D$S3�3��t$U�D$�D$������������Au������� ��}|  ���؋������� ��f|  ���؋��F��O�QP�R��O�Q��FP�R�N��j UPj j �?+ȋFQ�N�+�PWSQ���Da  ][��O�N�BPQ�PP��_�~(�ub�V,;V0tZ�D$P���D$  �?�D$    �D$     �|`  ����_  P���_  Pj j ���`  ���_  Pj j ���_  P����_  �F(���Q  9F$��   hh��L$(��S  hX��L$��S  �N(Q�T$xR�hV  �N$��P�D$(PQ�T$pR�QV  P�D$(P�L$lQ�aT  ��P�T$PR�ST  ��P�D$<P�ET  �N ��P�Z  �L$4�S  �L$D�S  �L$T�S  �L$d�S  �L$t�|S  �L$�sS  �L$$�jS  ^�Ā   � hD��L$�"S  h<��L$(�S  �V(�L$QR�D$\P�U  P�L$4Q�T$xR�S  ��P�D$|P�S  �N ��P��Y  �L$t��R  �L$d��R  �L$T��R  �L$$��R  �L$��R  ^�Ā   � �D$�T$�A�Q� ����������������D$V��L$�F$�D$���N(tc�F��t\��O�JPP�QH����t;W�~W��B  �T$�D$��j�Ή�F,�Y_  ��O�F�QPP�RP��_^� �L$Q�B  ��^� �D$�A0� ������VW���W  �N�����~D���  3��7�FH�FL�FP_����v0��^Ð���������V���   �D$t	V��h  ����^� ��V��N�����������V  ^Ð�����V��NP��t�q�����t�NP�u����NP��t�j��FP    ^Ð���������������AHÐ�������������V��h���L$�Q  �D$P��� X  �L$�'Q  jZjxj?h N  ���Z  ��u+h���L$��P  �L$Q�9a  ���L$��P  3�^���j�T$�D$R�FP���D$�����Z  ��u+h���L$�P  �L$Q��`  ���L$�P  3�^��ø   ^��Ð���������������ALÐ������������AL   Ð�������V���8����Ԗ��^Ð�������������V���   �D$t	V�[g  ����^� ���Ԗ�U������������O���   Vj ��L$j ����D$u)h���L$�O  �D$P�`  ���L$��O  ��   h(�h�   j�f  ����t�L$ �T$Q�L$RQ�VDR�������3����FPu)h��L$�IO  �D$P�_  ���L$�cO  �   ����R��u&h���L$�O  �D$P�{_  ���L$�/O  �Uj h�   h,  h,  h�  h�q j����T  ��u&h���L$��N  �L$Q�-_  ���L$��N  ��FH   �FH��u9�NP��t������t�NP�����NP��t�j��D$P�FP    �+K  ���FH^��� ��������������V���X���3��FT�F`� ���^Ð�����V���   �D$t	V�{e  ����^� ��� ��u��������V��jd��T  ����X  ^Ð�������������T$�D$��V��L$�V\�V`BW�FT�NX�~P�ωV`����j ����Z  ���pS  ��uUPh,  h�  h�  h�  h�q j���yS  ��u.h���L$�gM  �D$P��]  ���L$�M  _3�^��� _�   ^��� ������������V��FT���R  �NP��t�#������>  �NP��t�j��NT�FP    ��O���   j j ����D$�FT    u)h���L$��L  �L$Q�+]  ���L$��L  �   h(�h"  j ��c  ����t�V`�N\R�VXQ�L$RQ�VDR��������3����FPu&h��L$�]L  �D$P��\  ���L$�wL  �8����R��u&h���L$�,L  �D$P�\  ���L$�FL  ��FH   �FH��u9�NP��t�
�����t�NP�����NP��t�j��D$P�FP    �H  ��^��� ���������     Ð�������D$�T$�	P�D$R�T$PR������� ����������������	�9�������������	����V  �������	����V  ������h�Oj ��O��q  Ph�3j j �ĐP��O�ȐÃ�P��S3�V�t$\�L$(Q�D$,0   �D$0    �D$4�\$8�\$<�t$@�\$D�\$H�\$L�\$P�D$T���\$X��f��uhx��������^3�[��P� SVSSjdh�   SSh  � h��h��j��;ã�OuhX�������^3�[��P� P���;ã�Ouh(��o������_  h��P��;�uh���M������=  ��Oh��PR����uh���$������  ��OP�X�;ã�Ouh�����������   ��OPQ�ԑ��uhH���������   9��uh��������   UW��O�D$���D$���D$���D$���D$ ���D$$���D$(l��D$,P��|$�   �7V�}4  ����uVh8���������O��Mu�h��R4  ������_��O]��OSP�ԑ��OQ�ؑ��OR���^3�[��P� ���OÐ�����������OÐ�����������$ �����T  P�}���������   ��$X  ��$\  QR��$\  P�u���������   V3��L$Q�T$RVVVVVV��$x  P�L$|Q�D$<D   �t$@�t$D�t$H�t$hf�t$n�t$p�t$0�t$,�0���u1�8�Vh�   �T$`RVPVh   �`��D$XPh���i������L$�5ȐQ�֋T$R��^��T  Ð���������SVW�|$����1  ����Ǌ���:�u��t�P�^��:�u������u�3����������2  ���Ǌ���:�u��t�P�^��:�u������u�3���������l2  ����Ǌ���:�u��t�P�^��:�u������u�3���������02  ����Ǌ���:�u��t�P�^��:�u������u�3����������  �5��ht�օ���I��0  h\�օ���I��0  hD�օ���I��0  h,�օ���I��0  h�օ���I�|0  h�
�օ���I�h0  h�
�օ���I�T0  h�
�օ���I�@0  h�
�օ�� J�,0  h�
�օ��J�0  h�
�օ��J�0  hl
�օ��J��/  hT
�օ��J��/  h<
�օ��J��/  h$
�օ��J��/  h
�օ��J��/  h�	�օ�� J��/  h�	�օ��$J�x/  h�	�օ��(J�d/  h�	�օ��,J�P/  h�	�օ��0J�</  h|	�օ��4J�(/  hd	�օ��8J�/  hL	�օ��<J� /  h4	�օ��@J��.  h	�օ��DJ��.  h	�օ��HJ��.  h��օ��LJ��.  h��օ��PJ��.  h��օ��TJ��.  h��օ��XJ�t.  h��օ��\J�`.  hx�օ��`J�L.  h\�օ��dJ�F/  _^[þD�Ǌ���:�u��t�P�^��:�u������u�3��������u2�5��h,�օ��hJ��-  h�օ��lJ��.  _^[þ�Ǌ���:�u��t�P�^��:�u������u�3����������.  ���Ǌ���:�u��t�P�^��:�u������u�3���������`.  ���Ǌ���:�u��t�P�^��:�u������u�3����������   �5��h4��օ��pJ��,  h��օ��tJ��,  h���օ��xJ��,  h��օ��|J��,  h��օ���J��,  hl�օ���J��,  hP�օ���J��-  _^[þ8�Ǌ���:�u��t�P�^��:�u������u�3���������R-  � �Ǌ���:�u��t�P�^��:�u������u�3���������-  ��Ǌ���:�u��t�P�^��:�u������u�3����������,  ���Ǌ���:�u��t�P�^��:�u������u�3����������,  ���Ǌ���:�u��t�P�^��:�u������u�3���������b,  ���Ǌ���:�u��t�P�^��:�u������u�3��������uZ�5��h��օ���J�+  h|�օ���J��*  h`�օ���J��*  hD�օ���J��+  _^[þ,�Ǌ���:�u��t�P�^��:�u������u�3����������  �5��h�օ���J�l*  h�օ���J�X*  h��օ���J�D*  h��օ���J�0*  h��օ���J�*  h��օ���J�*  h��օ���J��)  h��օ���J��)  hx�օ���J��)  hd�օ���J��)  hP�օ���J��)  h<�օ���J��)  h$�օ���J�|)  h�օ���J�h)  h��օ���J�T)  h��օ���J�@)  h��օ���J�,)  h��օ���J�)  h��օ���J�)  h|�օ���J��(  hd�օ���J��(  hL�օ���J��(  h4�օ���J��(  h�օ���J��(  h�օ���J��(  h��օ�� K�x(  h��օ��K�d(  h��օ��K�P(  h��օ��K�<(  h��օ��K�((  ht�օ��K�(  h\�օ��K� (  hD�օ��K��'  h,�օ�� K��'  h�օ��$K��'  h��օ��(K��'  h��օ��,K��'  h��օ��0K��'  h��օ��4K�t'  h��օ��8K�`'  hx�օ��<K�L'  hd�օ��@K�8'  hP�օ��DK�$'  h4�օ��HK�'  h�օ��LK��&  h��օ��PK��&  h��օ��TK��&  h��օ��XK��&  h��օ��\K��&  h��օ��`K��&  h`�օ��dK��&  h@�օ��hK�p&  h �օ��lK�\&  h �օ��pK�H&  h� �օ��tK�4&  h� �օ��xK� &  h� �օ��|K�&  h� �օ���K��%  h� �օ���K��%  hl �օ���K��%  hL �օ���K��%  h< �օ���K��&  _^[þ( �Ǌ���:�u��t�P�^��:�u������u�3���������J  �5��h �օ���K�N%  h  �օ���K�:%  h���օ���K�&%  h���օ���K�%  h���օ���K��$  h���օ���K��$  h���օ���K��$  h���օ���K��$  ht��օ���K��$  h`��օ���K��$  hL��օ���K��$  h8��օ���K�r$  h$��օ���K�^$  h��օ���K�J$  h���օ���K�6$  h���օ���K�0%  _^[þ���Ǌ���:�u��t�P�^��:�u������u�3����������$  ����Ǌ���:�u��t�P�^��:�u������u�3����������$  ����Ǌ���:�u��t�P�^��:�u������u�3��������uh���������K�d$  _^[þ���Ǌ���:�u��t�P�^��:�u������u�3��������uhx��������K�$  _^[þd��Ǌ���:�u��t�P�^��:�u������u�3��������uhP��������K��#  _^[þ8��Ǌ���:�u��t�P�^��:�u������u�3���������|#  ���Ǌ���:�u��t�P�^��:�u������u�3��������u2�5��h��օ���K�"  h���օ���K�#  _^[þ���Ǌ���:�u��t�P�^��:�u������u�3����������"  ����Ǌ���:�u��t�P�^��:�u������u�3��������un�5��h���օ���K�v!  h���օ���K�b!  h���օ���K�N!  h���օ���K�:!  hl��օ���K�4"  _^[þP��Ǌ���:�u��t�P�^��:�u������u�3��������u2�5��h8��օ���K��   h ��օ�� L��!  _^[þ��Ǌ���:�u��t�P�^��:�u������u�3����������!  ����Ǌ���:�u��t�P�^��:�u������u�3��������un�5��h���օ��L�*   h���օ��L�   h���օ��L�   h���օ��L��  hx��օ��L��   _^[þ`��Ǌ���:�u��t�P�^��:�u������u�3��������u2�5��hH��օ��L��  h0��օ��L�~   _^[þ��Ǌ���:�u��t�P�^��:�u������u�3���������>   � ��Ǌ���:�u��t�P�^��:�u������u�3���������^  �5��h���օ�� L��  h���օ��$L��  h���օ��(L��  h���օ��,L��  h���օ��0L��  hp��օ��4L�v  hX��օ��8L�b  h@��օ��<L�N  h(��օ��@L�:  h��օ��DL�&  h���օ��HL�  h���օ��LL��  h���օ��PL��  h���օ��TL��  h���օ��XL��  h���օ��\L��  hd��օ��`L��  _^[þD��Ǌ���:�u��t�P�^��:�u������u�3���������h  �0��Ǌ���:�u��t�P�^��:�u������u�3���������,  ���Ǌ���:�u��t�P�^��:�u������u�3����������  ����Ǌ���:�u��t�P�^��:�u������u�3��������uh��������dL��  _^[þ���Ǌ���:�u��t�P�^��:�u������u�3���������`  ����Ǌ���:�u��t�P�^��:�u������u�3���������$  ����Ǌ���:�u��t�P�^��:�u������u�3����������  �x��Ǌ���:�u��t�P�^��:�u������u�3����������  �`��Ǌ���:�u��t�P�^��:�u������u�3���������p  �<��Ǌ���:�u��t�P�^��:�u������u�3���������4  �$��Ǌ���:�u��t�P�^��:�u������u�3����������  ���Ǌ���:�u��t�P�^��:�u������u�3����������   �5��h���օ��hL��  h���օ��lL��  h���օ��pL�l  h���օ��tL�X  h���օ��xL�D  h���օ��|L�>  _^[þx��Ǌ���:�u��t�P�^��:�u������u�3��������uhh��������L��  _^[þT��Ǌ���:�u��t�P�^��:�u������u�3����������   �5��h@��օ���L��  h,��օ���L�n  h��օ���L�Z  h ��օ���L�F  h���օ���L�2  h���օ���L�  h���օ���L�
  h���օ���L��  h���օ���L��  _^[þ���Ǌ���:�u��t�P�^��:�u������u�3��������uF�5��hp��օ���L��  h\��օ���L�x  h@��օ���L�r  _^[þ(��Ǌ���:�u��t�P�^��:�u������u�3���������2  ���Ǌ���:�u��t�P�^��:�u������u�3����������  ����Ǌ���:�u��t�P�^��:�u������u�3����������  ����Ǌ���:�u��t�P�^��:�u������u�3���������~  ����Ǌ���:�u��t�P�^��:�u������u�3���������B  ����Ǌ���:�u��t�P�^��:�u������u�3��������un�5��h���օ���L��  h���օ���L��  hh��օ���L��  hL��օ���L��  h,��օ���L��  _^[þ ��Ǌ���:�u��t�P�^��:�u������u�3����������   �5��h��օ���L�8  h���օ���L�$  h���օ���L�  h���օ���L��  h���օ���L��  h���օ���L��  h���օ���L��  _^[þ���Ǌ���:�u��t�P�^��:�u������u�3����������  ����Ǌ���:�u��t�P�^��:�u������u�3���������R  �p��Ǌ���:�u��t�P�^��:�u������u�3����������   �5��hT��օ���L��  h8��օ���L��  h��օ���L��  h���օ���L��  h���օ���L��  h���օ���L��  _^[þ���Ǌ���:�u��t�P�^��:�u������u�3����������  �5��h���օ���L�0  h���օ�� M�  ht��օ��M�  hd��օ��M��  hT��օ��M��  hD��օ��M��  h4��օ��M��  h$��օ��M��  h��օ��M��  h��օ�� M�|  h���օ��$M�h  h���օ��(M�T  h���օ��,M�@  h���օ��0M�,  h���օ��4M�  h���օ��8M�  h���օ��<M��  h���օ��@M��  h|��օ��DM��  hl��օ��HM��  hX��օ��LM��  h@��օ��PM��  h,��օ��TM�x  h��օ��XM�d  h ��օ��\M�P  h���օ��`M�<  h���օ��dM�(  h���օ��hM�  h���օ��lM�   h���օ��pM��  h���օ��tM��  hl��օ��xM��  hX��օ��|M��  hD��օ���M��  h0��օ���M��  h��օ���M�t  h��օ���M�`  h���օ���M�L  h���օ���M�8  h���օ���M�$  h���օ���M�  h���օ���M��  h���օ���M��  ht��օ���M��  h\��օ���M��  hD��օ���M��  _^[þ(��Ǌ���:�u��t�P�^��:�u������u�3���������z  ���Ǌ���:�u��t�P�^��:�u������u�3���������>  ���Ǌ���:�u��t�P�^��:�u������u�3����������   �5��h���օ���M��  h���օ���M��  h���օ���M��  h���օ���M��  h���օ���M��  h|��օ���M�v  h`��օ���M�p  _^[þD��Ǌ���:�u��t�P�^��:�u������u�3���������0  �,��Ǌ���:�u��t�P�^��:�u������u�3��������u2�5��h��օ���M��  h ��օ���M��  _^[þ���Ǌ���:�u��t�P�^��:�u������u�3��������u2�5��h���օ���M�f  h���օ���M�`  _^[þ���Ǌ���:�u��t�P�^��:�u������u�3��������u2�5��h���օ���M��  ht��օ���M��  _^[þX��Ǌ���:�u��t�P�^��:�u������u�3���������  �5��h@��օ���M��  h(��օ���M�z  h��օ���M�f  h���օ���M�R  h���օ���M�>  h���օ���M�*  h���օ�� N�  h���օ��N�  hx��օ��N��  hT��օ��N��  h0��օ��N��  h��օ��N��  h���օ��N��  _^[þ���Ǌ���:�u��t�P�^��:�u������u�3��������u2�5��h���օ��N�H  h���օ�� N�B  _^[þl��Ǌ���:�u��t�P�^��:�u������u�3��������uhT�������$N��  _^[þ<��Ǌ���:�u��t�P�^��:�u������u�3����������  ���Ǌ���:�u��t�P�^��:�u������u�3���������r  � ��Ǌ���:�u��t�P�^��:�u������u�3���������6  ����Ǌ���:�u��t�P�^��:�u������u�3����������  ����Ǌ���:�u��t�P�^��:�u������u�3����������  ����Ǌ���:�u��t�P�^��:�u������u�3����������  ����Ǌ���:�u��t�P�^��:�u������u�3���������F  ����Ǌ���:�u��t�P�^��:�u������u�3��������uZ�5��hh��օ��(N��	  hP��օ��,N��	  h<��օ��0N��	  h,��օ��4N��
  _^[þ��Ǌ���:�u��t�P�^��:�u������u�3���������x
  ����Ǌ���:�u��t�P�^��:�u������u�3����������  �5��h���օ��8N�	  h���օ��<N� 	  h���օ��@N��  h���օ��DN��  h���օ��HN��  h|��օ��LN��  h`��օ��PN��  hL��օ��TN��  h4��օ��XN�t  h��օ��\N�`  h��օ��`N�L  h���օ��dN�8  h���օ��hN�$  h���օ��lN�  h���օ��pN��  h���օ��tN��  h���օ��xN��  hh��օ��|N��  hP��օ���N��  h8��օ���N��  h��օ���N��  h ��օ���N�p  h���օ���N�\  h���օ���N�H  h���օ���N�4  h���օ���N�   h���օ���N�  h���օ���N��  hl��օ���N��  hX��օ���N��  hD��օ���N��  h0��օ���N��  h��օ���N��  h��օ���N��  h���օ���N�l  h���օ���N�X  h���օ���N�D  h���օ���N�0  h���օ���N�  h���օ���N�  h|��օ���N��  hh��օ���N��  hT��օ���N��  h@��օ���N��  h,��օ���N��  h��օ���N��  h��օ���N�|  h���օ���N�h  h���օ���N�T  h���օ���N�@  h���օ�� O�,  h���օ��O�  h|��օ��O�  hd��օ��O��  hL��օ��O��  h4��օ��O��  h��օ��O��  h��օ��O��  h���օ�� O��  h���օ��$O�x  h���օ��(O�d  h���օ��,O�P  h���օ��0O�J  _^[þt��Ǌ���:�u��t�P�^��:�u������u�3���������
  �\��Ǌ���:�u��t�P�^��:�u������u�3����������  �D��Ǌ���:�u��t�P�^��:�u������u�3����������  �0��Ǌ���:�u��t�P�^��:�u������u�3���������V  ���Ǌ���:�u��t�P�^��:�u������u�3���������  ���Ǌ���:�u��t�P�^��:�u������u�3����������  ����Ǌ���:�u��t�P�^��:�u������u�3��������uZ�5��h���օ��4O�~  h���օ��8O�j  h���օ��<O�V  h���օ��@O�P  _^[þ���Ǌ���:�u��t�P�^��:�u������u�3��������uhh�������DO��  _^[þ���Ǌ���:�u��t�P�^��:�u������u�3��������un�5��hT��օ��HO��  h@��օ��LO��  h(��օ��PO�p  h��օ��TO�\  h���օ��XO�V  _^[þ���Ǌ���:�u��t�P�^��:�u������u�3��������uF�5��h���օ��\O��   h���օ��`O��   h���օ��dO��  _^[þl��Ǌ���:�u��t�P�^��:�u������u�3��������u>�5��h���օ��hOtxhx��օ��lOthh`��օ��pO�b  _^[þD��Ǌ���:�u��t�P�^��:�u������u�3��������uh(�����tO���  _^3�[þ��Ǌ���:�u��t�P�^��:�u������u�3��������u$�5��h���օ��xOt�h���֣|O떾���Ǌ���:�u��t�P�^��:�u������u�3��������tt�P��Ǌ���:�u��t�P�^��:�u������u�3��������t<����Ǌ���:�u��t�P�^��:�u������u�3�������������_^�   [Ð�������O��SUVW�D$   �  h  �\������3������Ihh����D$�I3��������t�`�P�׋�����D$3����I�ٍD+P��P  �Ѓ��҉�Ouh�   h�h��P  ��j��O  ���3������+����������ȃ���O�|$�) ��O����D* 3����+��у�����=�O����O�ʃ�󤡄O��D( ��O��D) �D$��u_^]�   [���P�� ��O�����3��������I�҉t$��u��S�P  ������3������I;�v��SR�JK  ���Љ�O��uh�   h�h��O  ��j��yN  V� ��  �������   �}  ��   U�  �؊� ��OPU�T$(�   ����tU��������u_���3������+��у�����=�O�O�����ʃ����������+��у�����=�O����O�ʃ��t$�D$�D$U��u  P�?  ������G���V�_I  �D$��_^][��Ð������������SU�l$VW���3������AQ�N  �����3��������+������������ȃ����3�������+������у������O�ʃ��L�Ŋ��:u��t�P��:Vu������u�3��������uCh  �\���hHV�ZO  ��;��E  hDV�DO  ��;��/  _^]�   [þ4�Ŋ��:u��t�P��:Vu������u�3��������uCh  �\���hHV��N  ��;���   hDV��N  ��;���   h0�n���� �Ŋ��:u��t�P��:Vu������u�3��������uMh  �\���hHV�lN  ��;�t[hDV�ZN  ��;�tIh0V�HN  ��;�t7h������D$SP�,N  ����St�RG  ��_^]�   [��@G  ��_^]3�[Ð���D$���t�� t
��	t��
u�H@��u�Ð��������������D$���t�� t��	t��
t�H@��u�Ð��������������%��% ��%$��%��% ��%������������̡�O�H�!��������O�HV�t$�R�Q���    ^Ð���O�P�D$P�D$P�D$PQ�R��� �����������������O�P�D$P�D$P�D$PQ�R ��� �����������������O�P�D$P�D$P�D$PQ�R0��� �����������������O�P�D$P�D$P�D$P�D$PQ�R@��� ������������O�H�!��������O�HV�t$�R�Q���    ^Ð���O�P�D$P�D$P�D$P�D$P�D$P�D$PQ�R��� ��O�P�D$PQ�R��� �����������O�PQ�RYÐ���O�Hj��Q��Ð����������������O�T$�HR�QYÐ���������������OV��Hj�V���   ����^Ð�����T$��OV��HRV���   ����^� ��OV��Hj�V���   ��O�L$�Bj VQ���   ����^� ��������������O�PQ�RYÐ���O�PQ�R��á�O�P�D$PQ�Rh��� �����������O�P�D$PQ�Rt��� �����������O�P�D$PQ�Rl��� �����������O�P�D$PQ�Rp��� ����������T$��OV��HRV�Ql�����u3�^� ��O�QPV�R|��^� ���������VW�|$��W�r������u	�D$_^� ��O�HWV�QH��_^� ���������������VW�|$��W�2������u	�D$_^� ��O�HWV�QL��_^� ���������������VW�|$��W��������u	�D$_^� ��O�HWV�QD��_^� �����������������VW�|$��W�������u"�L$ �1�D$�Љ2�q�r�I_�J^��� ��O�BW�L$VQ�P`�Ћ2�D$$�ȉ1�r���q�R_�Q^��� ����VW�|$,��W�?������u�D$0�t$(P����  _��^��� ��O�QWV�RT���L$�D$,�b  �D$,��t
P�L$��  �D$,P�f  �t$,���L$Q���  �L$�  _��^��� ��VW�|$��W�������u�L$��D$��I_�H^��� ��O�BW�L$VQ�PX�Ћ
�D$ ����R_�P^��� ����O�P�D$P�D$PQ�R$��� ������O�P�D$P�D$PQ�R(��� ������O�P�D$P�D$PQ�R ��� ������O�P�D$P�D$PQ�R<��� ������O�P�D$P�D$PQ�R,��� ������O�P�D$P�D$PQ�R0��� ������O�P�D$P�D$PQ�R8��� ������O�P�D$P�D$PQ�R4��� ������O�P�D$P�D$PQ���   ��� ���O�P�D$PQ���   ��� ��������O�P�D$P�D$P�D$PQ���   ��� ��������������O�P�D$P�D$PQ���   ��� ���O�H$�a�������O�T$�H$R�QYÐ���������������OV��H$V�QD����^Ð�����������OV��H$V�QD�L$��O�B$QV�P����^� ��������OV��H$V�QD��O�L$�B$VQ�PL����^� ��������O�P$Q�RHYÐ���O�P$�D$P�D$P�D$PQ�R��� �����������������V��L$�a  ��O�H$V�Q�����D$t�T$R����  �D$P�  ���t$�L$Q���A  �L$�  ��^��� ����������������� V��L$�������O�H$V�Q �����D$t
P�L$�0   �T$R�   �t$,���D$P��������L$�������^�� � ���O�T$V��H$VR�QL����^� ����D$��VP�L$������O�D$,�Q$P�L$Q�R@�t$,���T$R���e����L$������^��Ð������O�P$�D$PQ�R<�����@� ����V�t$���t��O�Q$P�R���    ^Ð��������������O�H(�!��������O�H(V�t$�R�Q���    ^Ð���O�P(�D$P�D$P�D$P�D$P�D$P�D$PQ�R��� ��O�P(�D$P�D$P�D$PQ�R��� �����������������O�P(�D$P�D$PQ�R��� ������O�P(�D$PQ�R,��� �����������O�P(�D$PQ�R`��� �����������V�D$��P�D$    �D$    �������u^��� �D$��u(�L$�  �L$ P�Z  �L$�!  �   ^��� ��O�Qj j P��H  �����D$uj����=���3�^��� �L$j QP���������u�T$R�7  ��3�^��� �D$�L$j HPQ�L$,��  �T$R�  ���   ^��� ������������S�\$VW��j ���>  ��O�Hj Fj V��H  �����D$uj�������_^3�[� j VP���!  V���9   ��t�T$VR���H�����t�   �3��D$P�q  ��_��^[� ��������O�P(�D$PQ�R@��� �����������,V�t$4Vh�O�L$�  P�L$�������(����L$�o����L$�  ��^��,Ð���������������D$��O� Ð�����O�H@V�t$�R�QH���    ^Ð���O�PLQ�R ��á�O�PLQ�R$��á�O�PLQ�R8��Ã�0V��L$�!�����O�HL�T$Rj V�Q���L$�B����t$8Ph�  V�L$�~����L$�����L$�\�����^��0� �����V��L$�������O�HL�T$Rj V�Q��j h�  �L$�;����L$��������^��Ð����������V��L$�q�����O�HL�T$Rj V�Q���L$��  �t$$Ph�  V�L$�^����L$������^��� ��������������V��L$�����D$Ph�  �L$�^�����O�QL�D$Pj V�R���L$�^���^��� ���������O�H���   ����O�PL�D$P�D$P�D$PQ���   ��� ��������������O�PLQ���   ��Ð�������������L$�� ���������L$�T$�R�PÐ�T$�L$�R�T$R�PÐ������������T$�L$�R�T$R�T$R�T$R�PÐ��T$�D$Vh�}h�}h�}h�}R�Q�T$,R�T$,R�T$,R�T$,R�A�5�O�vLPQ���   ��,^� ��O�H�a�������O�T$�HR�QYÐ���������������OV��HV�Q`����^Ð�����������OV��HV�Q`��O�L$�BVQ�Pp����^� ��������OV��HV�Q`�L$��O�Bj j�QV�Pd����^� ����O�PQ�RlYÐ���O�P�D$PQ�Rp��� �����������O�T$V��HVR�Qp����^� ���V�t$���t��O�QP�R���    ^Ð��������������O�PQ�R��ËD$�L$��VPQ�L$��������"   �t$P��������L$�=�����^��Ð������D$V��P����P���;   ��^� �������O�P�D$P�D$P�D$PQ�R$��� �����������������O�P�D$P�D$PQ�R0��� ������V��L$�1�����O�T$$�H�D$ RPV�Q4�����D$t
P�L$�����L$Q������t$ ���T$R���	����L$�`�����^��� ���������O�P�D$PQ�R<��� �����������O�P�D$PQ�RP��� �����������O�P�D$P�D$P�D$PQ�RT��� �����������������O�T$V��H�D$R�T$PR�Q�����D$tP��������D$P�������������^� �����������L$������O�T$�HR�QD�����D$ t
P�L$�����D$ VP�����t$ ���L$Q��������L$�8�����^��Ð��VW�L$�2����D$$���|$ t%��O�Q4P�R����u6�L$����_3�^��Ë�O�B0W�P����u�L$�d���_3�^��Ë�L$Q�L$,Q���R$�L$���P������t��O�B0�L$QW���   ���L$����_��^��Ð�SVW�|$�������=ckhc��   ��   =TCAbatB=$'  t(=MicM�:  j hIicM��������WP���R_^[� �W���P_^�   [� j hdiem�������WP���R_^[� =INIbt=NIVb��   ����P_^[� �F��t_^�   [� ����F   �R_^[� ����P_^[� =ytsddtL=ndmct(=dmmc��   �Wj hidmc���)���P���S_^[� �Wj hidmc������P���S_^[� ����R _�F    ^3�[� =atnit$=cnysu"j hIicM��������WP���R_^[� ��  _^3�[� ��V���,���O�H0VhЁ��F���F    ��^Ð�����V���   �D$t	V��  ����^� ��V��F���,�t��O�Q0P�R���F    ^Ð��������O�P0�D$�IPQ���   ��� �����O�P0�Aj j j j j j j j j4P���   ��(Ð�������V��F��u^� ��O�Q0�L$ j j j j j Q�L$$j QjP���   ��O�B0�L$D�T$@Q�L$@R�T$@Q�L$<R�Vj QR���   ��D^� ������A��uË�O�Q0P�R��Ð�������A����Vu�t$P���  ��^��� �L$�Q�	�5�O�v0R�T$RQP�D$P���   �t$$��P���|  �L$�  ��^��� ������������O�P0�D$�IPQ�R ��� �������A��t(��O�Q0�L$j j j j j j Qj jP���   ��(� ���������������D$3҅���P�D$j BR�T$j PR�   � ��������������V��htniv�L$�����D$(Phulav�L$�)���hgnlfhtmrf�L$�����L$,Qhinim�L$�����T$0Rhixam�L$������D$4Phpets�L$������L$8Qhsirt�L$������D$$�T$RP�L$Q���d������m  �L$���R  �L$�y�����^��� ��V��hCITb�L$������D$(PhCITb�L$������L$,Qhsirt�L$�V����D$$�T$RP�L$Q�����������
  �L$����
  �L$������^��� �������������Q��u3�� �D$�H� V�5�O�v0Q�L$QPR�V8�L$3҃��ɋL$��^�� ���������������Q��u3�� �D$�H� V�5�O�v0Q�L$QPR�V8��^� ����������������Q��u3�� �D$�H� V�5�OW�|$Q�L$QP�|$�v0R�VD������t(�D$��t P�������L$��t���u���W�������_��^� �����Q�A��uY� ��O�D$     �Q0�L$ Q�L$j j Q�L$ Q�L$ Q�L$ j QjP���   �D$(��(Y� ��OV�t$�VW���H4R��D$�F    �~�H� ��O�R0Q�L$QVP�GP���   ��3Ʌ����F_^��� ���������D$��u��O� ��O�I�R0V�t$VP�D$PQ�RP��^� ����������������O�P0�Aj j j j j j j j j P���   ��(Ð��������   Ð����������   � ����������3�� T��H�H�HÐ�����������V���   �D$t	V�  ����^� ��V��FW3�;��T�u��O�V�H4R����~�~_^Ð����O�P4�AP�R��Ð��������������O�P4�AP�R��Ð��������������O�P4�AP�R��Ð��������������O�P4�D$�IP�D$P�D$P�D$PQ�R��� ���������O�P4�D$�IP�D$P�D$P�D$PQ�R��� ���������O�P4�D$�IPQ�R ��� ��������O�P4�D$�IPQ�R$��� ������VW�|$����!�����t��O�T$�H4�D$R�VPWR�QT��_^� �������������O�P4�D$(P�D$(P�D$(P�D$(�IP�D$(P�D$(P�D$(P�D$(P�D$(P�D$(PQ�RX��,�( �����������O�P4�AP�Rh��Ð��������������$V��F��tv�L$,��t(SW�x��O�X0���g���PW���   ��_[^��$� ���L���hARDb�L$�D$�D$    �����P�L$Q�N�T$R������L$��  �L$����^��$� ������V��h�  �����D$�L$�T$P�D$QRP���(���^� ����� �������������QSVW�|$���3�����=INIb��   ��   =SACb{t1=$'  t=MicM�I  _^��[Y� �W���P _�   ^��[Y� ��D$P�L$Q�Ή\$�\$�R��t��O�L$�B4�T$Q�NRQ�P��_�   ^��[Y� =ARDb��   USj���$���j j�ϋ�����j j�ϋ��
���j j�ωD$ ������P�D$PSU���R]_�   ^��[Y� ����R_�   ^��[Y� =NIVbYtB=NPIbt,=ISIbuP�>���h���P���@���P���W_�   ^��[Y� �W���P_^[Y� ����R_�   ^��[Y� =cnyst	_^��[Y� ShIicM���K����WP���R_^[Y� �����������V���x����|��F   ��^Ð������V���   �D$t	V�{  ����^� ���|����������VW�|$��������=cksat<=ckhct�D$PW������_^� ���F   ������t$_�F    �   ^� �F��t����R_^� _3�^� �����D$j0P�$   ��ËD$j$P�   �������@Ð���������O�T$�H�D$RP�QD��Ð��������O�H�T$�D$R�T$P�D$R�T$PRh4!  ���   ��á�O�T$�HR�QYÐ���������������O�H�ap�������O�T$�H�D$RP��,  ��Ð�����O�P���D$ P�D$P�D$PQ��D  �L$���#���ÐQ�D$���	�\$�A�$�\/  �\$�D$�$�L/  �t$��  ��� ����������W����������t
����\$���D$�G����G����t���\$�D$�@�������   �D$�@�������   �D$�������tS�D$�������tB�D$V�L  �D$���A  �ȋƙ����ҋ�u�t$�D$^�����G���__�؃���D$�D$�A/  �L$�T$�@��L$����At���t$��G�t$�__����    �G  �?_��Ð�������     �@  �?��D$V�������� ��$��-  ������F  zD������^� �����������qÐ������������     �@    Ë��L$�    �H� ���������������T$V���    �F    ��O���   j RV�Q����^� ���O���   Q�Yá�O���   Q�R8��Ð��������������O���   Q�R<YÐ����������������O���   Q�R@��Ð������������j�)   ����t�@��t�L$�T$Q�L$RQ�Ѓ��3�Ð���D$h�OPhD �  ��Ð�������Vj\�����������t�@\��tV�ЋD$��P���&   ��^� Vj`����������t�@`��tV�Ѓ�^�Vjd����������t�@d��t�L$QV�Ѓ�^� ����������   �����������3���O��O��OÐ�������������Vjp���&�������t�@p��t�L$QV�Ѓ�^� ��O^� j���������t	�@��t��3�Ð�����V�t$�> t!j���������t�@��tV�Ѓ��    ^Ð��Vj����������t�@��t�L$QV�Ѓ�^� 3�^� ���Vj,���v�������t�@,��t�L$�T$QRV�Ѓ�^� 3�^� ��������������Vj(���6�������t �@0��t�L$�T$Q�L$RQV�Ѓ�^� 3�^� �����������O���   �D$P�D$P�R� �������O���   �D$P�D$P�D$P�R� ��O�P �D$PQ�R��� �����������O�P Q�RYÐ�V�t$���t��O�QP�R���    ^Ð�������������D$�L$%�   S�؊���W�|$������f���ʃ��_[ËD$��s�   ��O�Qj j P��H  ��Ð����������D$��s�   ��O�Q�L$Q�L$QP��H  ��Ð����D$��t��O�QP�RYÐ����������V�t$ V�L$�����V�  ����t�L$Q�H �PL�t$�T$R��������L$�������^��Ð������   @� ���������   � ����������   U��$�   ��u��$�   �"���3�]�Ġ   �W3��`������D$��   SV��$�   P�L$(�a���h\�L$����P�L$D�I����t$Wj��L$,Q�T$LR��$�   P�������P��$�   Q������P�T$lR������P���A�����K��ۍL$\���O����L$x�F�����$�   �:����L$@�1����L$�X����L$$����^��[t0��$�   �L$��$�   UP��$�   Q��$�   RPQ�>   �����T$R�o�������$�   �D$    �������_]�Ġ   Ð���������������   V��$�   ��u
3�^���   �j �D$h�   P�S�����$�   ��$�   ��$�   h�   �L$T�L$Q�T$\��$�   �D$��$�   RPj�t$D�D$(0��D$lИ�D$p���D$t��D$x �������� ^���   Ð�����������`����������̋�`����������̋�`����������̋�`����������̋�� ��Ð���������Ð����������t�j�Ð�����D$��u��O�L$P�D$PQ�s�����Ð����������������3ɉ�H�H�H��   �����������V��F��Wu:���t��O�Q<P�R���    �~��t������W�e������F    _^Ð���������V�D$P���@�����P���   �L$���������^��Ð��V��F��W�|$u-h`j;j���������t
W���d����3����Fu_^� �F��t�3���_��^� ��O�H<W���3҅��_�F   ^��� �������������u��O�H�� ��O�J<�T$RP�Q��� ������   �   ��������O����������h��  YÐ�����O������������O�����������D$P��O�q���ø   � ��������3�� ������������ �������������� ���������������   V��$8  W���
�������$,  tj VW��������u	_^��   �j �D$h   P�������$P  ��$L  ��$@  Q��$H  RPQ�T$$R�+   ��$P  h   �D$,PQWj������4_^��   Ð�����D$�L$�T$V�t$P�D$Qj RPV�O  ��ǆ�   @�ǆ�   ��ǆ�   Мǆ�   ��ǆ�   �ǆ�    �ǆ�   �ǆ�    �ǆ�   0�ǆ�   ��ǆ�   ��^Ð�������������`\����������̋�`<����������̋�``����������̋�`@����������̋�`D����������̋�`H����������̋�`L����������̋�`P����������̋�`T����������̋�`X����������̋�`8����������̸   � ��������3�� ������������D$�L$�T$�H4�L$�P �T$��L$�@0��@8И�@<���@@��@D ��@H���@Lp��@P��@h ��@X0��@\@��@``��@dP��@T ��P0�H(�@,    Ë�`����������̋�` ����������̋�`$����������̋�`(����������̋�`,����������̋�`0����������̋�`4����������̋�`����������̋�`����������̡�O�PHjQ�Rd��Ð���������������� ���@    �V���   �D$t	V�[�������^� �������O�Px�AP�RYÐ����������OV��V�HxR�Q�D$����u	�   ^� ��O�Qx�L$Q�L$QP�D$P�3Ƀ������F^��� ��������������O�PXQ�R$��ø   � ��������3�� �����������3�� �������������   W3��������D$��   ��$�   SVP�L$$����h\�L$�����P�L$@�����t$Wj��L$(Q�T$HR��$�   P�-�����P��$�   Q�������P�T$hR�������P��������K��ۍL$X�������L$t������$�   �|����L$<�s����L$�����L$ �a���^��[t@��$�   �L$��$�   WP��$�   Q��$�   R��$�   P��$�   QRP�    �� ���L$Q��������_�Ġ   Ð�����   V��$8  W����������$,  tj VW�F�������u	_^��   �j �D$h   P������$T  ��$L  ��$P  Q��$D  R��$L  PQR�D$(P�3   ��$T  h   �L$0QRWj
�)�����8_^��   Ð�������������D$�L$�T$V�t$P�D$Q�L$RPQV�������ǆ�   @�ǆ�   ��ǆ�   М^Ð��������j�9   ����t+�@��t$�L$�T$Q�L$R�T$Q�L$R�T$QR�Ѓ��3�Ð����D$h�OPhD �|  ��Ð��������D$��Vu^Ët$�    �����u^É�@^Ð��������D$��t��T$�R�PÐ�����������D$��t�T$��R�T$R�PÐ������D$��t�T$��R�T$R�PÐ������D$��t�T$��R�T$R�PÐ������D$��t��T$�R�PÐ������������� ���@�@0��@`��@���@���@���@�Ð����������D$�T$jP�D$R��Q�L$PQ�q������ �����������3�Ð�������������D$�A � �������A Ð�������������V��NW���������u_�   ^��� �L$ �S�\$(UWSQ���P0�W�΋��R,��tWj htsem��������uEPhghcv��������u4Phrdem��������u#hﾭލL$�
����D$P���N����L$�U����L$(SQ������][_^��� ���������������D$��O�   � ����������������D$H����   �$�<��   á�S@����SuL�L$Q�������=L  }�����ËD$��u�����ÊV3���t��O+Ј�HF@��u�Ɔ�O ^�   ËT$�D$RP�$?���������H��>����Su
��>��������   Ã��ÍI ������5�����������������OÐ�����������O�HP�a@�������O�HPV�t$�R�QD���    ^Ð�V�t$��t���u9�D$jP�5�������u^Ë��E�����u^Å�t��p�T$3�;���I#�^Ð�������O�T$�HR���  ��Ð���������   ��  ��S�  ���ø��������������;��������U������}��f�E���f�E��m��}��m��E�U�����������̃��$�!  �   ��ÍT$�8!  R��<$tmf�<$t��   =  �?s-����������������=�S �Y!  �   ���V!  w8�D$��%�� D$u'��   ���t��������   ���� u�|$ u����- �   �=�S ��   �   ����  Z�����̃����$�T$�D$�   ��ÍT$�c   ��P��<$f�<$t�   ��  ��T$��  ���   �4   ��   �  ���   �L$���a  ����  ��u���=�S �T   ��   �   �=�S �7   ��   �)  ZÍT$��  �D$uA�3���   ���D$u����   �3��3�%�� D$uÍT$�  �D$��%  ����� =  �uT$u���u���t��Q���$�\$��q�"  ��Y�a���t����  �   �B����D$%�� D$������؋D$�  �t=�x   �l$���D$�   t�-0��t��   ���������0  ���)  ��%�� D$u���  ���  ���   ��������������- �   ���������ٱ ����u� �������ٛ���u������j��  Y�����������U��WV�u�M�}�����;�v;��x  ��   u������r)��$�ت�Ǻ   ��r����$���$����$�l�� �,�P�#ъ��F�G�F���G������r���$�ت�I #ъ��F���G������r���$�ت�#ъ�F��G��r���$�ت�I Ϫ���������������D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�ت��������E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$�p������$� ��I �Ǻ   ��r��+��$�x��$�p������Ы�F#шGN��O��r�����$�p��I �F#шG�F���G������r�����$�p���F#шG�F�G�F���G�������Z�������$�p��I $�,�4�<�D�L�T�g��D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�p������������E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_��V���   �D$tV�V���Y��^� VW�|$���ԗ�7��   @P�����Y�F��Yt
�7P��  YY�F   ��_^� VW�|$���ԗ�G���Ft%�w�   @P����Y�F��Yt�wP�y  YY��G�F��_^� �y �ԗt	�q����YËA��u�ܗ�V��j����5!  �vY��tV�J  Yj�!  Y^�V��������D$tV�g���Y��^� U��QSVW�E���E�d�    �d�    �E�]�c��m���_^[�� XY�$��XY�$��U��QQSVWd�    �E��E�:�j �u�u��u��  �E�@$��M�Ad�    �]��d�    _^[�� U���SVW��E�3�PPP�u��u�u�u�u�M!  �� �E_^[�E��]�U����E�e� �M�E�E�E��@�M��E�d�    �E썅����d�    �uQ�u�)  �ȋE�d�    ����U����Ej P�p�pj �u�p�u��   �� ]�U���4SVW�e� �E�Ư�E�E��E�E�E�E�E �E�e� �e� �e� �e� �E��e�m�d�    �E؍�����d�    �E�   �E�EЋE�EԍE�P�E�0�2)  �PhYY�e� �}� td�    ��]؉d�    �	�E�d�    �E�_^[��U��SVW��E�@��f��t�E�@$   jX�Mj�E�p�E�p�E�pj �u�E�p�u��  �� �E�x$ u�u�u������]�c�k �cjX_^[]�U��QSV�} W�}�w�_�Ɖu�E�|9���u��)  �MN��9L���};H~���u�E�M�E��u�} }ʋE��MF�1�M�;Gw;�v�~)  ��_^��[����U��SVWUj j hа�u�x�  ]_^[��]ËL$�A   �   t�D$�T$��   �SVW�D$Pj�hذd�5    d�%    �D$ �X�p���t.;t$$t(�4v���L$�H�|� uh  �D��@   �T���d�    ��_^[�3�d�    �yذu�Q�R9Qu�   �SQ�(�
SQ�(�M�K�C�kY[� U��� �EVWjY����}��E��E�E��E�P�u��u��u����_^�� U��V3�PPPPPPPP�U�I �
�tB�$��u����A�
�tF�$s���� ^��U��� �EV�E�E��E�E�B   P�E��u�E����P�)  ���M��x�E��  ��E�Pj �z(  YY��^�ËD$S��tJ�T$3ۊ\$��   t�
B2�tlHt.��   u��rW����ߋ�����_��t
�
B2�t>Hu�[Ã�r�
3˿���~����3σ��� �t��J�2�t#2�t��2�t2�t��_�B�[ÍB�_[ÍB�_[ÍB�_[áx�V��  �5�k��0  ��kY��k��+��;�s=R�0  ��P�5�k�  ����u3��,��k+�k��k������k�D$���k���  ��^��t$�y������Y��H�h�   ��  ��Y��kuj�  ��kY�  ��k��k�V�t$W����F@t�f �V�1  V�   V����1  ����_^�V�t$W����F�t4V�l3  V���3  �v�#2  ����}�����F��tP�  �f Y�f ��_^����������U��WVS�M�&�ً}��3����ˋ��u�F�3�:G�wtII�ы�[^_��U��V�u�1  �u�u�u�u�   �u���B1  ����^]�U��QSVW�}�}�]�υ��}��Mu3��   �uf�Ft�F�E��E   ��Mf�Ft*�F��t#;ȋ�r��W�6S�6  )})~>��ߋ}��K;Mr.�} ��t	3��u��+�PS�v�4  ����t6���t7)E��V� 3  ���Yt(��FC�M�E�} �v����E_^[�ÃN��N ��3�+E�u��V�:  ����u^�WV�t$�t$�t$�9  V���)0  ����_^�j@�t$�t$��������U��j�h�h�d�    Pd�%    ��SVW�u����   ��[��u;j	�  Y�e� V�=  Y�E��t	VP�=  YY�M���   �}� �Qj	��  YÃ�uSj	�^  Y�E�   �E�P�E�PV�J  ���E܅�tP�u��u���J  ���M���   �}� u�u�
j	�u  Y�Vj �5�[���M�d�    _^[��U��j�h0�h�d�    Pd�%    ��(SVW�]3�;�u�u�k  Y��  �u;�uS�����Y��  ��[���9  �}܃����   j	�  Y�}�S�<  Y�E�;���   ;5�[wLVSP�xD  ����t�]��8V�?  Y�E�;�t*�C�H�E�;�r��PS�u��4  S�8<  �E�SP�Y<  ��9}�uK;�uj^�u������uVW�5�[���E�;�t#�C�H�E�;�r��PS�u��3  S�u��	<  ���M���Z   9}�u";�uj^������uVSW�5�[���E܋E�;���  9=�T��  V�;N  Y��������  �u�]3�j	��  YÃ��G  ���w;�v������j^�u�}܃����   j	�-  Y�E�   �E�P�E�PS�H  �����}Ѕ���   ;52s\����SW�u��u��L  ����t�E�E��8S��H  Y�E܅�t*����E�;�r��P�u�u��2  W�u��u��jH  ���]�}� uSVj �5�[���E܅�t=����E�;�r��PS�u��N2  W�u��u��#H  ���VSj �5�[���E܃M���&   �E�;�uf9=�Tt^V��L  Y��������K�u�]j	�u  Y3��3����w;�uj^�����VSW�5�[��;�u9=�TtV�L  Y��u�3��M�d�    _^[�á���t��hD�h0���   h,�h ���   ���j j �t$�$   ���j j�t$�   ���jj j �   ���W�   j_9=(Tu�t$���P����|$ S�\$�=$T� Tu<��k��t"��kV�q�;�r���t�Ѓ�;5�ks�^hP�hH��C   YYh\�hT��2   YY��[t�   _��t$�=(T��_�j�  Y�j�  Y�V�t$;t$s���t�Ѓ���^�SV��WVj�*  V�WK  ���D$ P�t$ V�   VW����K  Vj�*  ��(��_^[��5�T�t$�   YYÃ|$�w"�t$�   ��Yu9D$t�t$��J  ��Yu�3��U��j�hH�h�d�    Pd�%    ��SVW��[��uC�u;5�[��   j	��  Y�e� V�,;  Y�E�M���   �E��tm�   j	�
  YÃ�uZ�E��t�p����j^�u;52w.j	�~  Y�E�   ����P�qE  Y�E�M���   �E��u-V��uj	�  YËE��ujX��$�Pj �5�[���M�d�    _^[������������̋L$WSV��|$��ti�q��tO���L$�F8�t��t�F8�t
��u�^[_3�ÊF8�u�~��a��t(���8�uĊA��t�f���8�t��3�^[_���#   �G�^[_Ë�^[_ÍB�[Í�$    �d$ 3��D$S�����T$��   t�
B8�tф�tQ��   u��W����V؋
����~����3���������3�3ƃ��� �u% �t�% u��   �u�^_[3�ËB�8�t6��t�8�t'��t���8�t��t�8�t��t��^_�B�[ÍB�^_[ÍB�^_[ÍB�^_[ËD$����   � �j��S�g4  ��Yt<��S3Ɋ�S%�   �-�S��S��S�����S��  ��u	�4  3��r�����k��M  �0T��H  �K  ��J  �r����,T�>3�;�u,9,T~��,T9$Tu�����SJ  ��  �4  ���uQ�J  YjX� U��S�]V�uW�}��u	�=,T �&��t��u"��k��t	WVS�Ѕ�tWVS�������u3��NWVS�+������Eu��u7WPS�������t��u&WVS������u!E�} t��k��tWVS�ЉE�E_^[]� �8T��t��u�=<Tu�N  �t$�8N  h�   ��YY�U��QQSV���  V�5��W  �EY�؋EYQf%�Qf=��$uU�:V  Y��Y~-��~��u#�ESQQ�$j�'O  ���pVS�FW  �EYY�b�E��SQQ�$�EQQ�$jj�=�U  �]��E��]YY���uVS�W  �E�YY�"�� u��E�SQQ�$�EQQ�$jj�	O  ��^[�������������̺���W  ���<W  �Ƀ=�St����c  �����z����h   h   �?g  YY�U����h��]��`��]��E��u��M��m��]��E������vjX��3���h������thp�P����tj �������V�t$�P�mh  ��eYt,F�=P5~�jP��g  YY���\5�A����uԊT5��F�����F��u�^ËD$�T5���t:�t�H@��u�@��t*���t��et��Et@���H�80t�8uH�@A�҈u�ËD$� �0����rjX�3��U��QQ�} �ut�E�P�pl  �EYY�M���M��H�ÍEP�l  �EYY�M���U���(�E�VP�E�P�EQQ� �$��l  �u�E�P�U�FP3��}�-��3Ʌ�����Q�]l  �E�j P�uV�u�	   �E��0^��U��S3�8]V�uW�}t3�9]��P3��>-���P�v  YY�>-��u�-�G9]~�P�H����T5�3�8]h�����MQ��	  9]YY��t�E�FA�80t<�^Ky���-A��d|��jd�^�� �Ù����A��
|��j
�^�� �Ù���� Y��_^[]�U���(�E�VP�E�P�EQQ� �$��k  �u�E�P�E��P3��}�-��EP�Ck  �E�j PV�u�	   �E��,^��U��SV�u�]W�FH�} t;Eu3Ƀ>-���ˋ�� 0�` �>-��u�-�{�F��jW�?  Y�0YG���} ~DjW�'  �T5Y��vGY��}+�} t�����9u|�u�uW��   �uj0W�"l  ��_��^[]�U���(SV�E�WP�E�P�EQQ� �$��j  �E�]�p�3��}�-��E���E�PSW�Bj  �E��H;������|&;�}"��t
�G��u� G��E�jPS�u���������E�jP�uS�u������_^[��U��}et2�}Et,�}fu�u�u�u�N�����]��u�u�u�u�4�����u�u�u�u������]�W�|$��tV�t$V�p  @PV�V�5�����^_���������������̀zuf��\���������?�f�?f��^���٭^�����剕l����ݽ`���ƅp��� ���a�����������$�����  ��؃��#�zuf��\���������?�f�?f��^���٭^�����剕l����ݽ`���ƅp��� �Ɋ�a�����ݽ`����Ɋ�a��������Ŋ�$׊���������$�����
�����  ��؃��#��   ������   ����������������۽b���ۭb�����i���@tƅp����ƅp�������۽b���ۭb�����i���@t	ƅp����ƅp������۽b���ۭb�����i���@t ��۽b���ۭb�����i���@t	ƅp����ƅp�����������- ��p��� ƅp���
��
�t���������U�����E��E�E��E�E��	U�����E��]��M�E�M�E�M�E�M�PQR�Qi  ���E�f�}t�m�����������������������������������ËT$��   ��f�T$�l$é   t�   �����   ËB%  �=  �t�ËB��
  ��D$�B�
�����D$�$�,$��
�    �BËD$%  �=  �tËD$�f�<$t�,$Z�f�$f=tf�� t���f�� t�   �����Z��,$ZÃ��$�D$��%  �����$�D$��%  �t==  �t_f�$f=t*f�� u!���f�� t�   ��t����Z��m���Z��,$Z��̘������������������   s��ܘ��Ę������������������   v��Ԙ�����ƅp����
�uK�����ƅp����2������;  ������a���t��=�St�����X  ��@u��
�t��������F  �t2��t�������������n��������-0ƅp����������ݽ`������a���Au����ƅp������-:�
�uS��������
�u�����~�����   ����
�u���u
�t���ƅp����-0��u�
�t��������=����������X��ݽ`������a���u���-0
�t���ƅp������������-0ƅp����
�u����-0������-N�ٛݽ`������a���Au�������ݽ`������a���������ݽ`�������������ٛ���u���b�����ٛ���t�   ø    ���   ��V��t��V���$���$��v�   ���f���t^��t������U��QQ�E�0��EV3�3����s���]��  ��  ��9Eu49UuW�E������we�E������rm��3�Ej^���   9Mu#9Uu�E������wB�E������s��9Eu19U��   �E�0����v��3�w�E�0����sg���e9Mue9Uu`�EQQ�$�X   �E�0�YY�����v��3��u���]�E�'�E�0����s��u��3����]�E���E���^��U��QQ�EQQ�$�(e  Y��YuI�EQQ�$�^I  �]��E��]YY���u,�E�58�QQ�]�E�$�5I  �]YY���uj�jX��3�������W�|$�j��$    ���L$W��   t�A��t;��   u�����~Ѓ��3�� �t�A���t#��t�  � t�   �t�͍y���y���y���y��L$��   t�A��td�G��   u���������~�Ѓ��3��� �t��t4��t'��  � t��   �t�ǉ�D$_�f��D$�G _�f��D$_È�D$_ËL$��   t�A��t@��   u�    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+��V�5��5����5����5����5���^�VW�=������t+���t#���t���t���tP���6�R���Y����P|��5����5����5����5���_^�U��EV�<�� �4��u>Wj������Y��uj����Yj������> YWu
���>������Yj�   Y_�6��^]�U��E�4����]����������̋T$�L$��   u<�:u.
�t&:au%
�t��:Au
�t:au����
�uҋ�3�Ð���@Ë���   t�B:u�A
�t���   t�f���:u�
�t�:au�
�t����U��V�uW� �9>t�?
  �E�@ft�~ to�} uij�V�u�u�  ���V�~ tP�8csm�u,9xv'�H�I��t�U$R�u �uV�u�u�uP�у� ��u �u�u$V�u�u�uP�
   �� jX_^]�U����E�e� �@����E�|�M;A|�	  SV�u�csm�W� �9�K  �~ub9~u]�~ uW��  �xl �&  ��  �pl��  �@pjV�E�E��Ha  Y��Yu�3	  9��   �~u9~u�~ u�	  9��   �~��   9~��   �}��E�P�E�PW�u �u��������؋E�;E���   9;|;{w�C�E�C���E�~d�F�@�x� ���E�~�v�7�u�=  ����u�M���9E���M�E�}� ��$�u��u$�u S�7�u�u�u�u�uV�  ��,�}��E����i����} t
jV�q  YY_^[�À} u �u$�u �u��u�u�u�uV�
   �� ���  U��QQVW�  �xh t!�u$�u �u�u�u�u�u���������us�}�E�P�E�PW�u �u����������E�;E�sO;>|C;~>�F�N����H��t�y u&j����u$�u Vj P�u�u�u�u�u�   ��,�E����_^��VW�|$�G��tJ�x �PtA�t$�N;�t��QR�Y���Y��Yu"�t�t�D$� �t�t	�t	�u3��jX_^�U��j�h�h�d�    Pd�%    ��SVW�e�]�s�u�};utU���~;w|�  �e� �G�D���th  SP�f  �M����u��/   YËe�M���}�]�u�G�4��u�릉s�M�d�    _^[�ËD$� �8csm�t3����  U��}  S�]VW�}t�u SW�u�  ���}, �uuW��u,������u$�6�u�uW�����Fh   �u(@�G�s�u�uW�u�   ��,��tWP�}���_^[]�U��j�h��h�d�    Pd�%    ��SVW�e�]�]ԃe� �u�F��E��+  �@l�E��   �@p�E��  �}�xl�
  �M�Hp�e� �E�   �u �uS�uV�������Eԃe� �M���:   �EԋM�d�    _^[���u��n   YËe�e� j��E�P�����YY3��ϋu�}�E؉F��  �M�Hl�  �M��Hp�?csm�u)�u#� �u�}� u�}� t�����PW��  YYËD$� �8csm�u�xu�x �u
�x ujX�3��U��j�h�h�d�    Pd�%    ��SVW�e�M�A���u  �x �k  �A���`  �U�|�e� �tD�uj�v�0\  YY���0  jW�:\  YY���  �F��M��QP�  YY��  �u�tR�]j�s��[  YY����   jW��[  YY����   �v�sW�������~��   �����   ��V뗃~ �]j�su:�[  YY����   jW�[  YY��t~�v��V�s��   YYPW�������f�R[  YY��tVjW�`[  YY��tH�v�n[  Y��t;�tj�FP�s�   YYP�vW�������FP�s�   YYP�vW��������  �M���M�d�    _^[��jXËe��g  U��j�h �h�d�    Pd�%    QQSVW�e�E��t�H�I��t�e� Q�p�`����M���M�d�    _^[��3�8E��Ëe��   �L$V�t$��Qƅ�|�42�I���^������U���SQ�E���E��EU�u�M�m��r���VW��_^��]�MU���   u�   Q�P���]Y[�� V������$�����`t:jtj�(Z  ��Y��Yt)V�5`� ���tV�4   Y���N�j�X^�3�^�������`���tP�(��`�ËD$�@P�7�@   �VW�8��5`���0�����u?jtj�Y  ��Y��Yt&V�5`� ���tV����Y���N���j�g���YW�,���_^á`�����   V�t$��uP�0�����tl�F$��tP����Y�F(��tP����Y�F0��tP�~���Y�F8��tP�p���Y�F@��tP�b���Y�FD��tP�T���Y�FP=�7tP�C���YV�<���Yj �5`� �^�U��j�h0�h�d�    Pd�%    QQSVW�e�3��u������9p`t�E�   �����P`�u��jXËe�e� �M���    �Y  U��j�hH�h�d�    Pd�%    QQSVW�e�e� �d��t�E�   ���jXËe�e� �M���    �I���V�t$��8csm�u�xu�x �u�&�����T��tP�W  ��Yt	V��T�3�^� h��4���T��5�T�4��U��SV�u�F�^����   �@��   �t�f ���   �N$���F�F�f �e $�f��Fu"���t���uS�[  ��YuV�K[  Yf�FWtg�F�>+��H��NI���N~WPS�2Y  ���E�6���t�ˋ��������Z������ 2�@ tjj S�X  ���F�M��j�E_WPS��X  ���E9}_t�N ��E%�   � �F���^[]�U���H  SVW�}3��G�ۉu�u�}��  �M�3���M��u�3�9U���  �� |��x�Ê�@����3����`������E���  �$���M���ỦU؉U��U�U��U��x  �Ã� t;��t-��tHHt���Y  �M��P  �M��G  �M��>  �M���5  �M��,  ��*u#�EP��  ��Y�E��  �M��؉E��  �E��ˍ��DA���U���  ��*u�EP�  ��Y�E���  �M����  ���ˍDAЉE��  ��It.��ht ��lt��w��  �M��  �M��  �M� �  �?6u�4uGG�M���}�l  �UЋ\5�U����DA�t�E�P�u��P�  ���G�}�E�P�u��P�f  ���%  �Ã�g�  ��e��   ��X��   �x  ��C��   HHtpHHtl����  f�E�0u�M��u����u�����EP�  f�E�Y�ȉM���  ��u	�l�M��E�   ����N����  f�8 ��  @@���E�   �� �M�@������;ʉ}���   �E�   ��   f�E�0u�M�f�E��EPt;�0  P������P�8X  ���E��}2�E�   �)��Zt2��	t�H��  �  ��  Y�������E�   �������E���  �EP�  ��Yt3�H��t,�E�t� ��M��E��E�   �  �e� �M�� �  �h�E�P�   u��gu�E�   �E�ũ��E�u��H��M��@��E���P������P�E�P���u�����   t�}� u������P��Y��gu��u������P��Y������-u�M��������}�W�����Y��  ��i��   ����   H��   HtQ�������HH��   ����  �E�'   �<+����  ��u	�h�M�����N��t�8 t@��+��  �E�   �E�   �E���E�   t]�E��E�0Q�E�   �E��H�E���E�   t;�M��5�EP�  �E� Yt	f�M�f���M��E�   �#  �M�@�E�
   �E��t�EP��  Y�A�E� t!�E�@�EPt��  Y����%�  Y�����E�@�EPt�  Y���  Y3��E�@t��|��s�؃� ���ڀM���������E��u�� �}� }	�E�   ��e�����u�e� �E��E��E��M������t;�E��RPWV�E��U��V  �uċ؃�0�u�WV�V  ��9����~]ԋE��M��뵍E�+E��E��E��E�t�M��90u��u�M�@�M��0�E�}� ��   �]���@t&��t�E�-���t�E�+�	��t�E� �E�   �u�+u�+u���u�E�P�uVj �  ���E�P�E��u�u�P�2  ����t��u�E�P�uVj0��   ���}� tA�}� ~;�E�]��x�f�CP�E�PC�YT  Y��Y~2�M�Q�uP�E�P��   ����O��u���E�P�u�u��u��   ���E�t�E�P�uVj �q   ���}�G�ۉ}�����E�_^[�Ú�p�������K���U��M�Ix��E�����Q�u����YY����Eu��]�� ]�VW�|$��O��~!�t$V�t$�t$�������>�t��O���_^�S�\$��KVW��~&�|$�t$�WF�t$P�u������?�t��K���_^[ËD$� � �@�ËD$� ��A��Q�ËD$� � f�@��U��j�hؙh�d�    Pd�%    ��SVW��[��uFj	����Y�e� �uV�  Y�E��t�v���	�u���u��M���	   �}� �U�u�j	����YÃ�uFj	�L���Y�E�   �E�P�E�P�u�  ���E؅�t�0���u���u��M���-   �}� u�uj �5�[�8����ƋM�d�    _^[�Ëu�j	�@���Yá�kVj��^u�   �;�}�ƣ�kjP�iM  Y��[��Yu!jV�5�k�PM  Y��[��Yuj�=���Y3ɸp��[��� ��=�|�3ɺ���������4��Z�������t��u�
��� A���|�^��H  �= T t�S  ËD$�p;�r=�w+�����P�����YÃ� P��ËD$��}��P�����YËD$�� P��ËD$�p;�r=�w+�����P����YÃ� P��ËD$��}��P�����YËD$�� P���V�t$;5�[s8�΋��������Z���D�tWV�U  V�(   V����U  ����_^��S  � 	   �
S  �  ���^�V�t$WV�U  ���Yt<��t��uj�U  j����T  Y;�YtV��T  YP�Ȑ��u
�8����3�V�TT  �ƃ���Y���Z���d� ��tW�R  Y����3�_^�V�t$�F��t�t�v����f�f��3�Y��F�F^�V�t$V�#   ��Yt���^��F@t�v�U  ��Y^��3�^�SV�t$3�W�F�ȃ���u7f�t1�F�>+���~&WP�v��L  ��;�u�F��t$��F��N ����F�f �_��^[�j�   Y�SVWj3�3������3�Y95�k~t��[����t_�@�tYPV������[YY���H���t0�|$uP�������YtC��|$ u��tP�������Yu���[�4�V����YYF;5�k|�j�����|$Y��t��_^[�V�t$�F����   �@��   �t
 �F�   f��Fu	V��M  Y��F��v�v�v�   ���F��to���tj�V�u7�NW���t�������<��Z�ɍ<��� 2�O_�ႀ��u�� �V�~   u�N��t��u�F   �H�F�A�^��������	F�f ���^�V�t$;5�[s@�΋��������Z���D�t%WV�{R  �t$�t$V�(   V����R  ����_^���O  � 	   ��O  �  ���^�U����e� �} S�]VW����  �E�ȃ����4����Z�<��Z��ƊH����  ��Ht�@<
t�M���S�E�   �D0
�E�j P��uR�40�<���u9�8�j^;�u�=O  � 	   �;O  �0���m�$  P�N  Y����  ��U�U��L0�D0����   ��t	�;
u�$���E�M��E�;��M���   �E� <��   <t�C�E�   I9Ms�E@�8
u�E�^�C�E�s�E�j P�E�E�jP��40�<���u
�8���uG�}� tA��D0Ht�E�<
t��C�D1�);]u�}�
u�
�jj��u��H  ���}�
t�C�M�9M�G������t0��@u�+]�]��E��3�_^[���U��WV�u�M�}�����;�v;��x  ��   u������r)��$����Ǻ   ��r����$���$����$���� �L�p�#ъ��F�G�F���G������r���$����I #ъ��F���G������r���$����#ъ�F��G��r���$����I �����������������D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$��������0��E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$��������$�@��I �Ǻ   ��r��+��$����$�����������F#шGN��O��r�����$����I �F#шG�F���G������r�����$�����F#шG�F�G�F���G�������Z�������$����I D�L�T�\�d�l�t����D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$��������������E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_��U��QQSV�5�UW�}3ۉ]��]��<at<rt<w�"  �  �3Ƀ���	  ��jZ�GG:���   ;���   ����Trt`��+tE��t6��tH��   9]���   �E�   �� �9]���   �E�   �����@u}��@���us���������΀   낸   ��uY��r�����btHHt.��t��u@���u;��@�S���9]�u.�E�   �������<���9]�u�E�   �� @  �%������t3������̀����h�  �uQ�u�M  �ȃ�;�}3���E��T�p�X��X�X�H_^[��SVWj3�3��m���3�9�kY��   ��[��;�t7�@�u!PV�S���YY��[���@�tPV����YYF;5�k|��_�<��Dj8������Y��[���[�;�t:�� P����[��� P����[�<;�t�O��_�_�_��_j����Y��_^[�V�t$j �& ��f�8MZu�H<��t��H��@�F^�U��,  ��P  ��h���SPǅh����   �H���t��x���u��l���rjX�  ������h�  Ph��D�����   3ۍ�����8�����t�<a|<z, �A8u퍅����jPh��~�������u�������I��d���h  PS�@�8�d�����d���t�<a|<z, �A8u퍅d���P������P����YY;�t>j,P�
���Y;�Yt0@��8t�9;u��A8u�j
SP�M  ����t��t��t�E�P�����}�Y���[��3�j 9D$h   ��P�ؐ����[t6��������[uh�  ��   Y�
��u�  ��u�5�[�L�3��jXá�[V��WufS3�9�[U�-�~@��[�=Ԑ�ph @  h   �6��h �  j �6���vj �5�[�Ճ�C;�[|��5�[j �5�[��][�'��u"�����F��th �  j P�Ԑ�6;�u��5�[�L�_^�h@  j �5�[������[uËL$�%�[ �%�[ j��[��[��[   Xá�[����[��;�s�T$+P��   r����3��U����MSV�u�AW�����+y����i�  ��D  �M��I���M���  �1�1�U�V��U��U����]u~��J��?vj?Z�K;KuL�� s�   �����L��!\�D�	u(�M!�!�J�   ���L��!���   �	u�M!Y�M��]��M��S�[M�Z�U�M��Z�R�S����J��?vj?Z�]����]���   +u��]���j?�uK^;�v��M��щM���J;�v��;�tc�M�q;qu@�� s�   �������!t�D�Lu&�M!1��K�   �����!���   �Lu�M!q�M�q�I�N�M�q�I�N�u��]�}� u;���   �M��\��щ^�N�q�N�q�N;Nu`�L�� �M���Ls%�} u�   �����M	�   �����D�D	�)�} u�J�   ���M	Y�J�   ��ꍄ��   	�E���D0��E����   ��[����   ��[�5Ԑ��H� �  h @  SQ�֋�[��[�   ���	P��[��[�@����    ��[�@�HC��[�H�yC u	�`���[�x�uiSj �p�֡�[�pj �5�[����[��[�����ȡ�[+ȍL�Q�HQP蒲���E����[;�[v�m��[��[�E�=�[��[_^[��U�����[��[SV��W�<��E�}��H����M���I�� }�����M���u��������3���u�E���[��;߉]s�K�;#M�#��u��;]��]r�;]�uy��;؉]s�K�;#M�#��u����;�uY;]�s�{ u���]��;]�u&��;؉]s�{ u����;�u�8  �؅ۉ]tS��  Y�K��C�8�u3��  ��[�C�����U�t����   �|�D#M�#��u7���   �pD#U�#u�e� �HD֋u�u���   �E�#U�����#9�t�U���3�i�  ��D  �M�L�D#�u����   j #M�_��|��G���M�T��
+M���M���N��?~j?^;��  �J;Jua�� }+�   �����M��|8�Ӊ]�#\�D�\�D�u8�]�M�!�1�O�   ���M��|8����   ��!��]�u�]�M�!K��]�J�z�}� �y�J�z�y��   �M�|���z�J�Q�J�Q�J;Jud�L�� �M})���} �Lu�   �����	;�   �����M�	|�D�/���} �Lu�N�   ���	{�M�����   �N�   ���	7�M���t�
�L���M��u�эN�
�L2��u��ɍy�>u;�[u�M�;�[u�%�[ �M���B_^[�á�[��[VW3�;�u0�D�P��P�5�[W�5�[��;�ta��[��[��[��[h�A  j���5�[�4���;ǉFt*jh    h   W���;ǉFu�vW�5�[��3���N��>�~��[�F����_^�U��Q�MSVW�q�A3ۅ�|��C����j?i�  Z��0D  �E��@�@��Ju��j��yh   h �  W�����u����   �� p  ;�w<�G�H�����  ����  �@��  ��������Hǀ�  �     �H�;�vǋE��O�  j_�H�A�J�H�A�d�D ����   �FC�������E�NCu	x�   �������!P��_^[��U����M�ESVW�}�׍p+Q�A�������i�  ��D  �M�O�I;�M�\9��|9��]��_  ���O  �;��E  �M���I��?�M�vj?Y�M��_;_uH�� s�   ���M��L��!\�D�	u+�M!�$���   ���M��L��!���   �	u�M!Y�O�_�Y�O��y�M+�M��}� ��   �}��M��O�L1���?vj?_�]���]�[�Y�]�Y�K�Y�K�Y;Yu\�L�� �M���Ls!�} u�   �����M	�D�D�   ����%�} u�O�   ���M	Y����   �O�   ���	�U�M��D2���L���U�F�B��D2��G  3��C  �:  �])u�N�K��\3��u�]��N�K���?vj?^�E���   �u���N��?vj?^�O;OuG�� s�   �����t��!\�D�u(�M!�!�N�   ���L��!���   �	u�M!Y�]�O�w�q�O�w�q�uu��u��N��?vj?^�M�|���{�K�Y�K�Y�K;Ku\�L�� �M���Ls!�} u�   �����M	9�D�D�   ����%�} u�N�   ���M	y����   �N�   ���	�E��D�jX_^[�Ã=�SUVWu���h    j �5�[�������  �-��jh    h  @ j �Ջ�����   j�   h   SW�Յ���   ��;�u�=� u���=� u�������F�5��F�0��  @ ���   �F�F�N�~�F3��   3҃���J#�JE��H����   |�Sj W�0  ���F�;�s���   ��G��G�   ��   �܋��'h �  j W�Ԑ���tVj �5�[��3�_^][�V�t$h �  j �v�Ԑ952u�F�2���t �F�Vj ���N�H�5�[��^Ã�^�U��QSV�5�W�~���   �e� ��   � �? �?�   u9��h @  Fh   P�Ԑ��t����T�F��t;�v�~�E��Mt��   ����}��}� �΋vt,�y�u&j�A Z�8�uB����   |��   uQ� ���Y;5�t
�} �P���_^[�ËD$��V��;Av;Ar�	;�t7��u1��   ���  ;�r �t$��t$��f�� �+��+�^���D�3�^ËD$�L$+H���D��L$��! �8�   �@�   u��T�=�T uj����Y�U��QQSV�52W�V�����   �~��   ��+ƃ������;��E�s:��];�|9_vSQP�  ����uu�E��_����      ;��E�r���]�F�N�~�E�;��M�s3�;�|9_vSP�u��j  ����u&�_�E�   ��;}�r���]�6;52t�C����52)�~�(  ������t� u�?;���   ��_�e� ���+�������w�;�u�}�}���E��8�t�E�j��h   PV�E����;���   j �u�V�F-  �U����ҋ�~0�F�U����   ��P�P���   ���A�      ���M�u։=2��   ;�s�9�t����;��#��G�E�F�_))F�L��   ��4�4�����t)�H�Y�T�2���   +ӉQ��)P��   �3�_^[��U��Q�M�USV�qW�9���   ;�}��ǉ]r!��;�s)Q�	�a �A��G��   ��> t�ƍ4;�sC���u0j�X^�; uCF��;�sN;E�u�q�)u9U��   �}������ƍ4;ur��q;�s~�;Esv���u@j�^X�; u%C@���;]s	+��q�	�a �q�1����6;�s)E9Ur4������맍;]s	+�A�	�a �A���Fk���+��3�_^[��U��Q�US�]V�
W�}�e� ��+G��;M�|�v�E+Ȉ�G�   �`se�E�4���   ;�rU�;�s
�8 u@��;�uB�E��;�w+;�v'���   ;�s3��38u@�< t��C�	�c �C�+M�E�   �E�_^[���VC20XC00U���SVWU��]�E�@   ��   �E��E�E��E��C��s�{���ta�v�|� tEVU�k�T�]^�]�t3x<�{S襪�����kVS�ڪ�����vj�D��]������C�T��{�v�4�롸    ��   �U�kj�S蚪����]�   ]_^[��]�U�L$�)�AP�AP�u�����]� ��T��t�t$�Ѕ�YtjX�3��V�t$�v�/0  ��Ytw���u3�����ucjX��Tf�FuR�<��T SW�<��T�   u S������Y�u�Fj�F�X�F�F��?�^�~�>�^f�NjX_[^�3�^Ã|$ Vt �t$�FtV�@����f�f �& �f Y^�U���HSVWh�  �
�����Y��uj����Y�5�Z��[    ���  ;�s�f ���f �F
��Z��$�  �ލE�P���f�}� ��   �E����   �8�X�;�E��   ;�|��9=�[}V��Zh�  �v�����Yt<��[ ����  ;�s�` ���` �@
���$���  ����9=�[|���=�[3���~L�E�����t8��t2�uQ�����t#�΋��������Z�����M��	���H�E�FC;�|�3ۋ�Z�ۃ<���4�uM���F�uj�X�
��H������P��������tW�����t%�   �>��u�N@���u
�N��N�C��|��5�[���_^[��SVW��Z���t7���  ;�s!�_�{� tS�����$�  ��$;�r��6蘬���& Y�����[|�_^[�S3�9�kVWu�<  �50T3��:�t<=tGV�'���Y�t���   P�α����Y;�5Tuj	�����Y�=0T8t9UW�������YE�?=t"U虱��;�Y�uj	蒵��YW�6�����Y��Y�8u�]�50T����Y�0T�_^��k   [�U��QQS3�9�kVWu��;  ��Th  VS�@���k�5T��8t���E�P�E�PSSW�M   �E��M���P���������;�uj����Y�E�P�E�P�E���PVW�   �E���H�5 T_^��S[��U��M�ESV�! �uW�}�    �E��t�7���}�8"uD�P@��"t)��t%�����Yt���t��F@���tՊ�F�����t�& F�8"uF@�C���t��F�@�����Yt���t��F@�� t	��t	��	ū�uH���t�f� �e �8 ��   ��� t��	u@��8 ��   ��t�7���}�U��E   3ۀ8\u@C���8"u,��u%3�9}t�x"�Pu����}�}3�9U�U���K��tC��t�\F�Ku���tJ�} u
�� t?��	t:�} t.��t�����Yt�F@���F������Yt@��@�X�����t�& F�������t�' �E_^[� ]�QQ��USU�-��VW3�3�3�;�u3�Ջ�;�t��U   �(�����;���   ��U   �   ����   ;�u�Ջ�;���   f9��t@@f9u�@@f9u�+Ƌ=����SS@SSPVSS�D$4�׋�;�t2U�f���;�Y�D$t#SSUP�t$$VSS�ׅ�u�t$軨��Y�\$�\$V������S��uL;�u�����;�t<8��t
@8u�@8u�+�@��U�������Y;�u3��UWV�!�����W������3�_^][YYá8T��t��u*�=<Tu!h�   �   ��UY��t��h�   �   Y�U���  �U3ɸH2;t��A=�2|�V����;�H2�  �8T����   ��u�=<T��   ���   ��   ��\���h  Pj �@���u��\���h��P�i���YY��\���WP��\����D���@Y��<v)��\���P�1�������\�����;j�h�W�'8  ����`���h؜P������`���WP������`���hԜP������L2��`���P����h  ��`���h��P�@7  ��,_�&�E��L2j P�6褾��YP�6j����P���^��U��=�: u)�u�EQQ�$QQ���$�EQQ�$�uj�  ��$]��=*  h��  � !   �u��  �EYY]�U���X�u �EP�u�6  ����u"�E�e��P�EP�E �u�uP�E�P�]   ���u��  �=�: Yu,��t(�u �EQQ�$QQ���$�EQQ�$�uP��  ��$��P�h  �$��  �u �F  �EYY��U��M3�SV�A�MWj�A�M[�A�M��t�E�E�  �	X��t�E�E�  ��H��t�E�E�  ��H��t�E�E�  ��H��t�E�E�  ��H�u�Ej��P��#˃�����_�H��E�ыP������ʉH��E�ыP������ʉH��E�ыP��#σ��ʉH��E�ыP��#˃��ʉH�'  ��t�M�I�t�M�I�t�M�I�t�M	y� t�E	X��   #�t4=   t=   t;�u(�E�� �E������
�E����ˉ��E� ���   #�t =   t;�u"�E� ���E�������E�������E�M���  ����� ��ʉ�E	X �E�H ���ωH �E� �E�X�E	XP�E�HP���ϋ}�HP�E��X@�%  �EPSj �u����E�@t�&��@t�&��@t�&��@t�&�Xt�&ߋ��������� t%ItIt	Iu�N����������������!������� tItIu!��#ʀ���#ʀ���@@�_^[]�U����ESW����j�[t�]tS�  Y�����  �t�Etj�s  Y����  ����   �E��   j�Q  Y�   �M#���   ��   tX��   t(;���   �M��0���3���w���]��E��n�M��0����v��3���3���]��E��F�M��0����v��3���3���]��E���M��0���3���w���]��E�������   ���   �E��   V3��t��E� �]��E��0������   �E�E�PQQ�$�I  �E����]� ���������}	����]��T�E��0����s���3ҊE���f�E�����;�}+��]�t��u���m�]�t�M���m�Hu��t�E����]��E�E�����^tj�  Y����Et�E tj �  Y���3���_[����U��� �u�   ��Y�E�tU�EV�E�E�E�E�u�E��Eh��  �u(�E�E �u��E��E$�E��'  �E�P�U  ����uV�$   Y�E�^��h��  �u(��  �u�   �E ���ËD$��t~���$$  � "   ��$  � !   �3ɸ�2�;T$t��A=�3|�3�Ë��2ÊD$� tj��tj��tj��tjX��������U��QQ�E���]��E���U��QQ�E�M�E�  f����]����f�E��E���U��3ҁ}  �u	9Uuj�<�}  ��u	9Uuj�*�M��  #�f;�uj�f���u�E�� u9UtjX]�3�]�U��QQ�E�0�V���u��3��]��   3�f�E�ue�E�� u9MtW�E�0��������sjX�3��Eu�e�E�t�M�eN��f�e��;�t�M��EQQQ�$������]����'�EQQQ�$������E���]���f%������  �E�E��0^��U��Q��}��E���U��Q�}����E���U��Q��}��E��#E��#M�ȉM�m�E���U��QQ�M��t
�-�3�]���t����-�3�]�������t
�-�3�]����t	�������؛�� t���]��������������U���0���S�ٽ\�����=�: t�׭����8����   [����ݕz������U���U���0���S�ٽ\����=�: t�3�����8�����8�����Z   [��ݕz�����U���0���S�u�u�  ���u�u�  ���ٽ\�����8���ƅq����<����   [�À�8�����=�S uLݕ0�����p���
�t<�t@<�t<
�t0����r����   f��\���f�� u���f�� tǅr���   �z٭\�����f��6���f%�f�tf=�t0�ǅr���   �؝�����������ȝ����s4���,ǅr���   �Н�����������������v���VW��l���C��v�����8���u��u��z������{t�u�}����]���r�����\���SP��l����C��P�  ��_^�E��$���U���0���S�u�u�   ���ٽ\�����8�����j�������[��U����Sf�Ef��f%�f=�uf���f�]��E�]���E��]��m���E[���������l$�l$�D$���   5   �   t��������3 u��ËD$%�  tg=�  t`�|$�D$?  %��  �D$ �l$ �D$%�  ��t� 4��� 4���l$����4���4���l$��ËD$D$u��ËD$%�  u��|$�D$?  %��  �D$ �l$ �D$%�  t=�  t2�D$�s*��D$�r �������4�|$�l$�ɛ�l$������l$��Ã�,��?�$�N4����,Ã�,�����,Ã�,�����,�����,�����,�����,��|$���<$�|$ �����l$ �Ƀ�,Ã�,��<$�|$�����l$�Ƀ�,Ã�,����|$���<$�|$ �^����l$ ��,��<$�|$�J�����,��|$�<$�:����l$��,��|$�<$�&�����,��|$�����<$�|$ �������l$ �ʃ�,Ã�,��<$���|$��������l$�ʃ�,Ã�,����|$�����<$�|$ ��������l$ ��,��<$���|$�����Ƀ�,��|$���<$�������l$��,��|$���<$�����Ƀ�,��|$�����<$�|$ �j������l$ �˃�,Ã�,��<$���|$�K������l$�˃�,Ã�,����|$�����<$�|$ �$������l$ ��,��<$���|$�����ʃ�,��|$���<$��������l$��,��|$���<$������ʃ�,��|$�����<$�|$ ��������l$ �̃�,Ã�,��<$���|$�������l$�̃�,Ã�,����|$�����<$�|$ �������l$ ��,��<$���|$�h����˃�,��|$���<$�T������l$��,��|$���<$�<����˃�,��|$�����<$�|$ �"������l$ �̓�,Ã�,��<$���|$�������l$�̓�,Ã�,����|$�����<$�|$ ��������l$ ��,��<$���|$������̃�,��|$���<$�������l$��,��|$���<$�����̃�,��|$�����<$�|$ �~������l$ �΃�,Ã�,��<$���|$�_������l$�΃�,Ã�,����|$�����<$�|$ �8������l$ ��,��<$���|$� ����̓�,��|$���<$�������l$��,��|$���<$������̓�,��|$�����<$�|$ ��������l$ �σ�,Ã�,��<$���|$�������l$�σ�,Ã�,����|$�����<$�|$ �������l$ ��,��<$���|$�|����΃�,��|$���<$�h������l$��,��|$���<$�P����΃�,Ã�,�<$�|$�;�����,Ã�,�|$�<$�(�����,�P�D$%  �=  �t3��% 8  t�D$����X� �Ƀ��<$�D$�����,$�Ƀ�X� �t$X� P�D$%  �=  �t3��% 8  t�D$�k���X� �Ƀ��<$�D$�V����,$�Ƀ�X� �t$X� P��% 8  t�D$�/���X� �Ƀ��<$�D$�����,$�Ƀ�X� P��% 8  t�D$�����X� �Ƀ��<$�D$������,$�Ƀ�X� P�D$%  �=  �t3��% 8  t�D$�����X� �Ƀ��<$�D$�����,$�Ƀ�X� �|$X� P�D$%  �=  �t3��% 8  t�D$�~���X� �Ƀ��<$�D$�i����,$�Ƀ�X� �|$X� P��% 8  t�D$�B���X� �Ƀ��<$�D$�-����,$�Ƀ�X� P��% 8  t�D$����X� �Ƀ��<$�D$������,$�Ƀ�X� P��,�<$�|$������,X�P��,�|$�<$�������,X�PSQ�D$5   �   ��  ������4 �p  �D$%  �=  ��\  �D$.%  ��M  =  ��B  �D$,��6  �D$��*  �D$%�  ��?�\$0���  +�w^�D$%�  ��
�\$0���  +���   �l$(�D$�\$0���  ��+؃���+ˋ؁� �  ˉL$�l$�D$�����|$(�����   u�l$�|$�|$4�D$4?  �D$8�l$8�D$%�  �\$0���  +؃�?�� ���ˋD$�\$0���  % �  ؉\$�l$���l$(������%   u�����<4�Ƀ�u�\$0�|$(���l$�-D4�����l$(�l$4�� �  t���
�l$�l$(����   tV�|$<��   t�|$4�D$4   �D$8�l$8�,4�l$4�D$<�����l$��% C  ���4$�d$��  	D$�$$��Y[X�R��0�|$�<$3ҋD$�  �t
�������0Z��,$�l$�$D$ty���|$�,$�Ƀ��|$$�D$$?  �D$(�l$(�D$ %�  =�  w���$4�|$�$4�<$� �|$$�D$$   �D$(�l$(���$4�<$�l$$�T�����0Z�����0Z�PSQ�D$5   �   ��  ������4 �p  �D$%  �=  ��\  �D$.%  ��M  =  ��B  �D$,��6  �D$��*  �D$%�  ��?�\$0���  +�w^�D$%�  ��
�\$0���  +���   �l$(�D$�\$0���  ��+؃���+ˋ؁� �  ˉL$�l$�D$�����|$(�����   u�l$�|$�|$4�D$4?  �D$8�l$8�D$%�  �\$0���  +؃�?�� ���ˋD$�\$0���  % �  ؉\$�l$���l$(������%   u�����<4�Ƀ�u�\$0�|$(���l$�-D4�����l$(�l$4�� �  t���
�l$�l$(����   tV�|$<��   t�|$4�D$4   �D$8�l$8�,4�l$4�D$<�����l$��% C  ���4$�d$��  	D$�$$��Y[X�R��0�|$�<$�    �D$�  �t
�������0Z��,$�l$�$D$ty���|$�,$�Ƀ��|$$�D$$?  �D$(�l$(�D$ %�  =�  w���$4�|$�$4�<$� �|$$�D$$   �D$(�l$(���$4�<$�l$$�Q�����0Z�����0Z�������@����������U��QV��}��u��:   ���E��#��E#E�V�   Y�EY�m��^�ËD$%����P�t$����YY�S�\$3�U��WtjX��t��t��t�� t��t   ��V�Ѿ   �   #ֽ   t��   t��   t;�u������#�^t;�u   �   _]��[t   �S�\$3�V��tjX��t��t��t��t ��   t�˺   #ʾ   t��   t;�t	;�u���������ˁ�   t��   u���^��   [t���U��Q�E�H��   w�\5�A�R��V�5\5�����DV�^t�e� �M��E�j�	�e� �E�jX�M
jj j QP�E�Pj��  ����u���E
#E��S3�9Vu�D$��A|Y��ZT�� [�V�`XWV���9\X�=��tV��j�֤��Yj[�t$�   ��Y�D$t
j����Y�V�׋D$_^[�U��Q�=V SVWu�E��A��   ��Z��   �� �   �]�   j;�^}%95P5~VS�����YY�
�\5�X#ƅ�u���e�\5�������DJ�t�e
 j�E�]	X�	�e	 �]��Vj �M�jQP�EPW�5V�&  �� ��t�;�u�E���E��M����_^[�ËD$Vj �Y��j���D$���Y�D$+ʃ�����҅�uF��}���8 uF����|�jX^�3�^ËD$SVWj �\$�Y�����D$����<�WjYjX+���P�7�2(  ��Nx�<���tWj�7�(  ��N����}�_^[�U��QQ�ESVW�x�j Y�e� �_j ��^���j�ȋÙ���E^j�M����E+�Z����t!CS�u����Y��YuW�u�N���Y�E�Y�E�������jY!�E�@;�}�U+ȍ<�3��E�_^[�ËD$�L$Vj+�Z�0�4��Ju�^�W�|$3����_ËD$3Ƀ8 uA����|�jX�3��U����ESVWj �}[�������E�   ���E�E����e ����+��֋��#ΉM�����E��E��˃����M��Eu܋}�j[��jY��;�|�U��+Ƌ���E�$ K��y�_^[��U����ESVW�H
�ف� �  �M�H�M�H� �}���  ���?  �M���������E�u&�E�3�P������Y��   �E�P�����YjX��   �E�P�E�P�����w�E�P��������tC�G��+O;�}�E�P����Y�<;�?+Ë��E�P�E�P�v����E�VP�����w�E�P������G@P�E�P������ 3��|���;|(�E�P�V����w�M���E�P�m����w��7j�R����w�w�e��E�P��I���YY3�jY+O���M��Ɂ�   ��u��@u�M�U��q��
�� u�M�1_^[��hh7�t$�t$�������h�7�t$�t$�l������U���3�PPPP�u�EP�E�P�&  �u�E�P������$��U���3�PPPP�u�EP�E�P�q&  �u�E�P������$��U��US�]V�u�JW�~�0�ۋ�~�]3ۊ��t��A�j0Z�@�Mu�U�  ��|�95|H�89u� 0��� �>1u�B�W�~���@PWV�Ez����_^[]�U���(V�EWP�E�P�G   Y�E�Y�u�Pj j������f��*  �u�}�F�Eډ�E؉F�E�PW�-����� �~��_^��U��Q�USVWf�B��  ��% �  ��#ωE�B��پ   �%�� �ۉu�t;�t�� <  �(��  �!3�;�u;�u�E�X�f�X�K��<  �]�������ȋEM����H���u�ɋ���ٍ��X����  ���ߋM�f�H_^[������������̋T$�L$��tG3��D$W����r-�ك�t+шGIu������������ʃ���t��t�GJu��D$_ËD$�j賎��Y�U���X�ESV�u��WH�Mt+Ht$HtHtHtHHtHunj��   �bj�
j�j�j[�~QWS��������uA�E��t��t��t�e����M��F����]Ѓ��M��NWQP�ESP�E�P������h��  �u������>YYt�=�: uV�l9  ��Yu�6�����Y_^[��U��E��  ��#�f;�u,�EQQ�$�c���YHYtHtHtjX]�j��j���   ]�% �  f�ҋ�u�E�� u�} t�����$��   ]��E�0������u���$���@]����$   ]�Vj^�t$�t$�����t3���^�Vj^�t$�t$�����t3���^�Vj^�t$�����t3���^�U��j�h�h�d�    Pd�%    ��SVW�u�u�u�u���w3�;�uj^������u�3ۉ]������   ��[��uA�}�;=�[w|j	�ڛ��Y�]�W�3���Y�E��M���   9]�t^�u��H3ۋuj	����YÃ�uA;52w9j	藛��Y�E�   ����P����Y�E��M���L   9]�tVS�u�������9]�u>Vj�5�[���E�9]�u'9�TtV�����Y���0����3ۋuj	腛��YËE��M�d�    _^[��j
����j�   YYj�r���V�t$;5�[s@�΋��������Z���D�t%WV�  �t$�t$V�(   V���^  ����_^��  � 	   �~  �  ���^�V�t$WV�  ���Yu�V  � 	   �-�t$j �t$P��������u�8��3���tP�  Y�����΃����Ƌ��Z���d���D���_^�V�t$;5�[s@�΋��������Z���D�t%WV�=  �t$�t$V�(   V���  ����_^��  � 	   �  �  ���^�U���  SVW3�9}�}��}�u3��f  �E�����Z�E���4�����D0 tjW�u����������@���   �E9}�E��}��   �������M�+M;Ms)�M��E��	��
u�E�� @�@�ȍ�����+ʁ�   |̋�������+��E�j P������WP��40�����tC�E�E�;�|�E�+E;Er�3��E�;���   9}tbj^9uuL�  � 	   �  �0�A�8��E�ǍM�WQ�u�u�0�����t�E�}�E���8��E��u��  Y����,��D0@t�E�8������!  �    �  �8��+E�_^[����Th   �̄��Y�L$���At�I�A   ��I�A�A�A   �A�a �ËD$;�[r3�Ëȃ��������Z�D���@�U��SV�`XWV����=��3�9\XtV��j蘗��Yj[�u�u�   Y�E��Yt
j�ڗ��Y�V�׋E_^[]�U��E��u]Ã=V uf�Mf��� w9j�X]ÍM�e Qj �5P5P�EjPh   �5V�����t�} t��  � *   ���]���SV�D$�u�L$�D$3���؋D$����A�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$vN3ҋ�^[� ��������S�D$�u�L$�D$3���D$���3��P�ȋ\$�T$�D$���������u�����d$��d$�r;T$wr;D$v+D$T$+D$T$���؃� [� SWj3�����Yj_9=�k~]V��[�������tA�@�tP��z�����YtC��|)��[��� P����[�4��|����[Y�$ G;=�k|�^j����Y��_[�V�v   �L$3���08;t"��F=�9|��r"��$w�B   �    ^��5   ��48^�Á��   r���   w�   �    ^��   �    ^���������
������QQSUVWj�������3�Y�\$�\$��Z�u ����   ���  ;�st�FuD�~ u#j�͔���~ Yu�FP���Fj����Y�^S���FtS���\$�E ��$�  륃���+E j$Y�����|$���um�\$�D$ ��C���[�\$�^����N��  V������Yt>��[ ���Z���  �;�s�` ���` �@
���$�������W�O  Yj�]���Y��_^][YYËL$V;�[WsU�����<��Z�����4�����<0�u6�=<TS�\$u�� tItIuSj��Sj��Sj��|���03�[��c���� 	   �a����  ���_^ËL$V;�[WsX�����<��Z�����4������@t7�8�t2�=<Tu3�+�tItIuPj��Pj��Pj��|���0�3�������� 	   ������  ���_^ËD$;�[s�ȃ��������Z�D���t� ������ 	   �����  ���ËD$S�ȃ���VW�4��Z���Z�<�����~ u#j胒���~ Yu�FP���Fj�ɒ��Y��D8P��_^[ËD$�ȃ��������Z�D�P���S�\$;�[VWsr�����<��Z�Ã��4�����D0tRS�J����Y�D0t)S�����YP�x���u
�8����3���t�����0����� 	   ���S�b���Y�������� 	   ���_^[�U����MS3�V���W�E�   �]�t	�]��E���e� �E�   � �  ��u��@u9$Vt�M��j��^#�+�tHtH��   �E�   ���E�   @��E�   ��E��t&�� t��0t
��@ut�u���E�   ��E�   ��]�   �   #ʿ   ;�1t*;�t&;�t��   tM��   u+�E�   �L�E�   �C�u��>��   t/��   t;�t#�q����    �o��������  �E�   ��E�   �E��   ��t��S��#M���uj^�@t
��   �M���t�� t��   �
�t��   �����؃��;�u������    ������  ���*  j V�u��E�P�u��u��u�t���;�u�8�P�<���Y����   V�����u	V�Ȑ�؃�u�M�@�	��u�M�VS������Y��Y�M��<��Z�À����M�4�����eH�L0ux���ts�Etmjj�S�����������E�u�.����8�   tKS�����Y����X�e �EjPS�.�������u�}u�u�S��  Y���Yt�j j S�m��������t��} u�Et��L0 �D0��S����Y��_^[��j �t$�t$�t$�   ���U���S�e� VW�}��w�u��=P5~��jP� ���YY��\5�ÊA����t�F�Ѐ�-�u�u�M���+u�F�u��E����  ����  ��$�w  j��Yu$��0t	�E
   �2�<xt<Xt	�E   ��M9Mu��0u�<xt<Xu�^FF�u����3��u�  �E�=P5��~jV�C���YY��\5�p����t�˃�0�2�=P5~WV����YY��\5f�p#ǅ�tJ��P�  Y�ȃ�7;Ms6�u��M;u�ru���3��u;�v�M�	�u�u��E��E���d����E�M��]�u��t�E�E��e� �K�����u�u>��t	�}�   �w	��u,9u�v'������E� "   t�M����E$�����ƉE���t�E���Et�E��؉E��E���E��t�83�_^[��������Q=   �L$r��   -   �=   s�+ȋą���@P�U���SVWj�q����u�  ��Y;dXY�]u3��p  ���V  3Ҹ�99tt��0B=�:|�E�PS�p�j^;��!  j@�%�Z Y3���Y9u�󫪉dX��   �}� ��   �M�����   �A���;���   ���Y@��e� j@Y3���Y�4R�������9�; ��t,�Q��t%���;�w�U����9��Y@;�v�AA�9 u��E����}�r��E�|X   P�dX��   ���9�pX��Y��Z��RAA�y� �G����ƀ��Y@=�   r�S�   Y��Z�5|X��%|X 3��pX�����=�U t�   �   �������j�=���Y��_^[�ËD$�%�U ���u��U   �%h����u��U   �%l����u�V��U   ËD$-�  t"��t��tHt3�ø  ø  ø  ø  �Wj@Y3���Y�3��pX�dX�|X��Z���_�U���  �E�VP�5dX�p����  3��   ������@;�r�E�ƅ���� ��t7SW�U��
��;�w+ȍ�����A�    �����˃��BB�B���u�_[j �������5�Z�5dXP������VPj�L  j �������5dXVP������VPV�5�Z��  j �������5dXVP������VPh   �5�Z�  ��\3�������f���t���Y���������X���t���Y �������〠�X @AA;�r��I3��   ��Ar��Zw���Y�Ȁ� ���X���ar��zw���Y �Ȁ� �����X @;�r�^�Ã=�k uj�����Y��k   �S3�9�UVWuBh8��d���;�tg�5�h,�W�օ���UtPh�W��h�W��U�֣�U��U��t�Ћ؅�t��U��tS�Ћ��t$�t$�t$S��U_^[�3������̋L$W��tzVS�ًt$��   �|$u��uo�!�F�GIt%��t)��   u����uQ��t�F�G��t/Ku�D$[^_���   t�GI��   ��   u����ul�GKu�[^�D$_É��It�����~�Ѓ��3��� �tބ�t,��t��  � t��   �uƉ�����  �����   ��3҉��3�It
3����Iu���u��D$[^_�U����E�e� HSVHWtgHHtF��tA��t<��t*��tHt����F  ��U��U�B��U��U�5��U��U�(萐�����vP�u�  ��Y��Y����U��Uj�E�   �n����uY��u�}� ��   S趆��Y��   3�;�u9M�tj螆��Yj�q���E��t
��t��u�VT���U��NTuI�VX�FX�   �U��u7�8�8�;�}(�I���VP���d� �8�=8A�;�|����}� tj����Y�}u�vXj��YY��u�Ӄ}Yt�}u�E��}�FTu�E�FX3�_^[�ËT$�$8V�t$9rW��t�<I�<���;�s9pu�I��;�s9pt3�_^�U��j�hP�h�d�    Pd�%    ��SVW�e��U3�;�u>�E�Pj^VhH�V�X���t����E�PVhD�VS�\�����   jX��U��u$�E;�u�V�u�u�u�uP�\��   ����   9]u�V�ESS�u�u�E �����@P�u�̐�E�;�tc�]��< �ǃ�$������e��u�WSV��������jXËe�3�3��M��;�t)�u�V�u�uj�u�̐;�t�uPV�u�X��3��e̋M�d�    _^[��U���   SV�u3�;��(  ���  j�҃���\XY9`Xt
j�А��;�Wt$9]t�uV��  YY��  �v�4��;��  �}�E�   ;��]��  �?L�  �C�  �_�  h��W�  ��Y;�Y��   �3ۋ�+ǉE���   �>;��   �E   ��;��E�PW�3�h������u�3�����9E�Yt�E�����;~�Fh��V��e����Y��Yu�>;u[�}/W��x���VP�������=x��� ��x���P�u��   ����t�E��? t.G�? t(h��W�  ��Y��Y�:���3�j�ׂ��Y3��   �} ��   3��   SS��x���SPW�m  ����;�tw��;��;�t/�7��x���P諂��Y��Yt��x���PS�d   Y��Yu!E���E��C���;~�3�9}�t�Y  �5�;���i��Y�=�;�9}�j����6  ��j�'���Y�\X��_�3�^[��U���   SVW�}�E�WP�E�P��\���P�u�  ������   ��\���P�f���@P�n��Y�E��Y��   �4�� V��j���;�E��E��EDV�E�P�E�P�����V�E���\���P�u������;j�E���E�P�u��ݝ���E�� ��u�V��u�V���;��t#�E�u���;��g���E�Y��E��V3���}�:t	�u��g��Y���;_^[�á�;SUVWj��]uhQ  �*m��Y��;�  �5�;���W�5�;j�5�;�  ��;����h���5�;�M~���v���3谀������t3��6��W�v�j�5�;�J  �����;|�_^��][u��;��5�;�g���%�; ��;Y�U���   SV�u3�;�W��   �>Cu28Vu-�E�M P;�� Ctf�f�Qf�Q�M;���   ���   �,;VW����Y��Ytt��:VS����Y��Ytb��x���VP�   Y��Yu��x���P��x���h�UP�  ����u3��i��U��U��x���PW�F  �> YYtV�WS�}��YY�} tjh�U�u�՛�����} tjh�U�u轛����W�u��|��Y��Y_^[��W�|$��~V�t$�v���t$�|��YOYu�^_�U��SVW�}h�   j W�-����u�����t<.u�~ �Ft�ǀ   PW�g|��YY3��   �e h��V�_a��Y��Ytj�} �0�<0u��@}Y��.tTPV�u�4�}u��@}B��_t=P�EV��@��}u-��t��,u$P�EV�   P���������,t���t��E�w녃��_^[]�V�t$V�t$��{���~@ �F@YYtPh��j�t$����������    ���   ^tPh��j�t$��������U��j�h��h�d�    Pd�%    ��SVW�e�3�9= VuFWWj[ShH��   VW�P���t� V�"WWShD�VW�T����"  � V   9}~�u�u�  YY�E� V��u�u�u�u�u�u�u�T���   ����   9} u�V�E WW�u�u�E$�����@P�u �̐�؉]�;���   �}����$�������e�ĉE܃M���jXËe�3��}܃M���]�9}�tfS�u��u�uj�u �̐��tMWWS�u��u�u�P����u�;�t2�Et@9}��   ;u�u�uS�u��u�u�P�����   3��eȋM�d�    _^[���E�   �6��$������e�܉]��M���jXËe�3�3ۃM���u�;�t�VS�u��u��u�u�P���t�9}WWuWW��u�uVSh   �u �����;��q������l����T$�D$��V�J�t�8 t@��I��u�8 ^u+D$Ë�ËT$V�t$3��2;�r;�sjX�T$^�
�V�t$W�|$V�7�6���������t�FPj�0��������t�F�FP�w�0��������t�F�FP�w�0������_^ËD$VW�0�x����0�4?���H�׉p�����_�H^ËD$VW�P�H�������ΉH��������_�P�^�U����ES�]3�;�V�E�N@  ��S�SvQW�E��}�S��p���S�j����E�PS����S�Z����E�e� �e� � �E��E�PS��������E�Mu�3�_9Su(�K�����C�����������E���  �s��Ӿ �  �suS������E���  Y��f�E�^f�C
[��U���\SVW�}�E�j�E�3�Z�E؉U�E��E��E܉E��EԉEЉE�E��E�}��� t��	t
��
t��uG��j^�G���w  �$��Y��1|��9j�  :T5uj�F  �Ã�+tHHt����  �   j�E� �  X맃e� jX란�1�U�|��9~�:T5��   ��+t1��-t,��0tR��C��  ��E~��c�{  ��e�r  j��  Oj��  ��1|	��9�V���:T5�Y�����0��  �������U�9P5~��VP����YYjZ��\5�ÊA#ƅ�t�}�s�E��E���0�E���E��G�:T5ug��������}� �U��U�u��0u�M��G��9P5~��VP�E���YYjZ��\5�ÊA#ƅ�t�}�s�E��E���0�E��M���G빀�+�
�����-���������9P5�U�~��VP�����YYjZ��\5�ÊA#ƅ���   ���W�O���1�M|��9~D�Ã�+ttHHtd���  j�e�U���0u�G����1��   ��9��   �
��1|��9	j	XO������0uD���}  t*�ÍO���+�MtHH��   �M��jX����jX����j
OX��
��   �o����}�   �E�   3��=P5~��jP�����YY��\5�ÊA����t�ˍ��tAЁ�P  �G뾾Q  �u�=P5~��jP����YY��\5�ÊA����t�G��O����E�}� �8��   jX9E�v�}�|�E��E��E�H�E���E�}� ��   H�8 u�M��E���E�P�E��u�P�j����E�3Ƀ�9M�}��E�9M�uE9M�u+E=P  ~0�E�   �]�u�E�U�}� t`3۸�  �   �3��E�   �^=����}	�E�   ���uP�E�P�  �U��]uƋEʃ��3�3�3�3��3�3�3�3��E�   ��}� t3�3�3�3��E�   �ME�_�q�Yf�A
�E�^f�[�æU�ULVvV�VHW~W�W�W,XX�WU����ES�]V�Ⱦ�  �� �  #�f��W�E���E���E���E���E���E���E���E���E���E���E���E�?�E�   ��t�C-��C �}f��u��u9}uf�# �C �C�C0��  f;�uz�   �f� ;�u�} t��   @uh��Ff��t��   �u�} u.h���;�u#�} uh؞�CP��q��Y�CY�e� �n  hО�CP��q��Y�CY���ϋ���i�M  ��f�e� j�Nf�U�k�M�}�����E���E�����P�E�P�  ��f�}��?r�E�FP�E�P�j  YY�Ef�3t�}�����������}��~j_�u����?  f�e� �E   �E�P�]����MYu��}�ށ��   ~�E�P�n���NYu�O�C�ɉE~P�M�u��}���E�P������E�P�����EP�E�P�����E�P������E��M�e� ��0�E�M�u��E�H�HH��5�K|0;�r�89u� 0H��;�s@f�� *�,�C���d �E�_^[��;�r�80uH��;�s�f�# �C �C�0�c jX��U��  �s���SV3�jV�u���������;ÉE���   jV�u�d�����;���   W�}+���~u�   ������SVP�p���h �  �u�p  ���E;���}��P������P�u����������t+���~���r����8u�_����    ����u�u�  YY�H}Fj �u�u������u�`�����P�L��������N;�u�����    �8����
����8j �u��u��������_���^[��S3�9Vu�D$��a|Y��zT�� [�V�`XWV���9\X�=��tV��j��p��Yj[�t$�   ��Y�D$t
j�q��Y�V�׋D$_^[�U��Q�=V Su�E��a��   ��z��   �� �   �]��   }(�=P5~jS�����YY��\5�X����u���k�\5�������DJ�t�e
 �E�]	j�	�e	 �]jX�M�jj jQP�EPh   �5V�n����� ��t���u�E���E��M����[�Ã=V VtZh�   j�m�����Y��YujX^�V�h   ��YtV�  V�V��YY���5(V�5xC�  �5(V�V��Y�5(VY�)�5(V�xC�C�f  �5(V�oV���%(V YY3�^�U��QQ�bV�dVV�u���E��M�u����"  S�NWQj1Pj[S�  ���FPj2�u�S�  ��FPj3�u�S��  ��FPj4�u�S��  ��@��FPj5�u�S��  ��FPj6�u�S�  Vj7�u��S�  ��F Pj*�u�S�  ��@��F$Pj+�u�S�  ��F(Pj,�u�S�v  ��F,Pj-�u�S�e  ��F0Pj.�u�S�T  ��@��F4Pj/�u�S�@  ��FPj0�u�S�/  ��F8PjD�u�S�  ��F<PjE�u�S�  ��@��F@PjF�u�S��  ��FDPjG�u�S��  ��FHPjH�u�S��  ��FLPjI�u�S��  ��@��FPPjJ�u�S�  ��FTPjK�u�S�  ��FXPjL�u�S�  ��F\PjM�u�S�  ��@��F`PjN�u�S�k  ��FdPjO�u�S�Z  ��FhPj8�u�S�I  ��FlPj9�u�S�8  ��@��FpPj:�u�S�$  ��FtPj;�u�S�  ��FxPj<�u�S�  ��F|Pj=�u�S��  ��@����   Pj>�u�S��  ����   Pj?�u�S��  ����   Pj@�u�S�  ����   PjA�u�S�  ��@����   PjB�u�S�  ����   PjC�u�S�s  ����   Pj(�u�S�_  ����   Pj)�u�S�K  ��@����   Pj�u�S�4  ����   Pj �u�S�   �ƨ   �Vh  �u�S�	  ��0�_[^��V�t$����  �v��R���v��R���v��R���v��R���v��R���v��R���6��R���v ��R���v$��R���v(�R���v,�R���v0�R���v4�R���v�R���v8�R���v<�R����@�v@�}R���vD�uR���vH�mR���vL�eR���vP�]R���vT�UR���vX�MR���v\�ER���v`�=R���vd�5R���vh�-R���vl�%R���vp�R���vt�R���vx�R���v|�R����@���   ��Q�����   ��Q�����   ��Q�����   ��Q�����   ��Q�����   ��Q�����   �Q�����   �Q�����   �Q�����   �Q�����   �Q����,^�S3�9VUW�=^V��   Vh,VjWj]U�E  h0VjWU���5  h4VjWU��%  �54V��k  ��4;�^t>�5,V�Q���50V�Q���54V�Q�����,V�0V�4V����4  �x� =@t#P��P���x�p��P���x�p�P�����x�,V��x�0V�H�x�4V�H�x� � �-X5�T5�   �5,V�iP���50V�^P���54V�SP��j�,V�0V�4V��U���x����x� ;��1���h��P��f��j�U���x���A�x�@;�����j��qU��Y�x�A�x�@;��������x� � �X5   �T53�_][Ã=V Vtvj0j�,�����Y��YujX^�V�   ��YtV��  V�xO��YY��x� ��x�@�F�x�@�F�58V�5x�  �58V�9O��Y�58VY�G�x�58V��H�H�L�@�P�xH�q  �58V��N���%8V YY3�^�V�t$W�=XV��u����  �FSPjWj�  �؍FPjWj�  ؍FPjWj�  ؍FPjWj�w  ��@؍FPjWj�d  �v��   �F PjPWj�L  ؍F$PjQWj�<  ؍F(PjWj �,  ��D؍F)PjWj �  ؍F*PjTWj �	  ؍F+PjUWj ��  ؍F,PjVWj ��  ��@؍F-PjWWj ��  ؍F.PjRWj ��  ��/�VjSWj �  ��0�[_^ËL$���tV<0|<9,0�A���u�^�<;u���P�p��ƀ8 u���V�t$��tC�F=�St9P�rM���v�jM���v�bM���v�ZM���v�RM���v �JM���v$�BM����^�U���$S3�9V�]��]���  9VVWu#�PVhVh  PS��  ������  �  V�rR����V�}��gR��h  �E��ZR��V�E��QR����;��E��t  9]��k  9]��b  ;��Z  3��   �M��@;�|��E�P�5V�p����0  �}��&  �E܃��P5~,8]�t'�E�:�t�H���;��U��A���@@8X�u�S�GSSPV�u�j����������   �M�f�3�f�AA@;�|��E�SS�xWV�u�j�  ������   �E�f��=P5~68]�t1�E�:�t(�p���;��M��Lqf� �F�AA;�~�@@8X�uҋE��=`5���\5�<V;�tP�K��Y�E�<V�@V;�tP�hK��Y�E��@V�u��WK���u��OK��Y��Y_^�L�u��?K���u��7K��YYj[���5<V�f5�\5�`5�K���5@V�K��Y�<VY�@V3�[��3����U��V3�PPPPPPPP�U�I �
�tB�$��u�
�t
F�$s�F��� ^��S3�9�VVWu�  ��t�@���V�
��V�r�t$;���   �5xV8thxVj@hpA�*  ���F@;ã|Vt8th|Vjh�@�  �|V���xV��V;�t8t;�t8t�5  ��  �;�t8t�  ��s  9�V��   �ƀ   V�u  ��Y;���   ��P�D�����   j�5hV�H���ts�D$;�tf�hVf�f��Vf�Hf�x�t$;�tEj@Vh  �5hV��V��t2�F@j@Ph  �5�V��V��t�ƀ   j
VW�2  ��jX�3�_^[�U��SVW3�9]jX|C��t?�EÙ+��E���4��<��E�0�  Y��Yu
�M���9�}N�u��^;]~�_^[]��5xV�`���5|V�����@�tV�`����Y����%hV @�=tV Y�lVt�pV   ��5xV�X  Y�pVjh�m�<���V��t	��t�u�%�V �U���xSVW�u��  Y���E�jxP�lV���f%�  PV��V���  �E�P�5|V�  Y������Y�  ��   �E�jxP�tV���#��PV��V����   �E�P�5xV�I  Y��Yuf��V�5�V�5hV�m��Vud�pV��t:P�E�P�5xV��  ����u#�5xV��V�5�V�;_��;pVYu#���VuV�K  ��Yt��V�5�V��V�   #�;���   �E�jxP�tV���#��PV��V��u�%�V jX�   �E�P�5xV�m  Y��Yu1��V3�9=tVuW9=pVtO�5xV�^��;pVYu;j�+3�9=tVuB�pV;�t9P�E�P�5xV��  ����u"WV�  Y��Yt��V9=hVu�5hV��V������_^[�� �5xV�^����Y���@�tVt�pV   ��5xV��  Y�pVjh�o�<���Vu�%�V �U���xV�u�  Y���E�jxP�tV���f%�  PV��V��u!�VjX�w�E�P�5xV�0
  Y��Yu9tVu:j�*�=tV u@�pV��t7P�E�P�5xV��
  ����u PV�  Y��Yt��V�5�V�5hV��V������^�� �5|V�]����Y���j@h�p�lV�<���Vu�%�V �U���xV�u�  Y���E�jxP�lV���f%�  PV��V��u!�VjX�@�E�P�5|V�<	  Y��YuV�   ��Yt��V�5�V�5hV��V������^�� f��V�,���V�hV�U��QQV�u��t1�> t,ht�V�]��Y��Ythp�V�]��Y��Yu(�E�jPj��E�jPh  �5�V��V��t
�u�V�[
  Y^�ø�@f�L$f;t@@=�@|�jX�3��U���x�E�jxP�E%�  j��P��V��t5�E�P�Q  9EYt*�} t$V�5xV�r  �5xV���e[��Y;�Y^u3���jX��U���   ��l���ǅl����   P�H���t��|���ujX��3���U��SVWj3�_�7�]�+�����k�,�� <9Mt(9Ms�x���p;�~�S�u�u�u�@�_^[]� �MIt[IItM��t>��t/���  tItIIu�k�,$<�<k�,��<�1k�,��<�&k�,<�k�,<�k�,<�k�,<���x������o����u�K�QPV�Y������d� jX�a����T$3��
B��t+��a|
��f������A|��F�������������ËT$3��
B��A|��Z~
��a|��z@���U���$S�]V�uf�K
3�W�E�E܉E��E�f�F
����  3�#�#ʁ� �  f=���U��  f�����  f������  f���?w3��:f������u�E�Vu3�9Fu9u�o  3�f;�u�E�Su9Cu9u�F�F��k  �E��E��E��E   �E���} ~IƍK�E��E�M�E�E��M�� �	���M����QP�1���������t�E�f� �E��m��M�uȃE��E��M�} ��E�  f�} ~%�E�u�E�P������E��  Yf�} �f�} 9�E��  f�} }+�E��E���E�t�E�E�P�����KYu�}� t�M�f�}� �w�E�%�� = � u5�}��u,�e� �}��u�e� f�}���u�Ef�E� ��f�E���E���EދEf=�sf�M��f��M��N�M�Nf�F
�f����f ��   ��� ���& �~_^[��U���S�0D3Ƀ�`9Mtc}�E��E�؉E��`9Mu�Ef�9MtAVW�E��T�}��;�t'�@f�<� ��4�r�}�����M��u�V�u�r���YY3�9Mu�_^[�ËD$V�ȃ������ �  ���Z�T��L���%�   9t$u����|$ @  u�ɀ����
f% ��^�������    ���^�U���   �}SVW��   3ۍE�Sh�   P�}��u�]�u��  ����;�uM�8���zu^SSS�u�u�  ����;�tGV�9D����Y;�t:SVW�E   �u�u�  ����;�tV�D��Y;ËM�u9]tW�q>��Y���_^[��VWP�=�����9]ttW�R>��Y�k�} u�j ��VjV�u�u�  ����t��}�' �=P5�~��jP�_���YY��\5�ÊA����t��
���,0FF����V|�3��p���U��j�h��h�d�    Pd�%    ��SVW�e衔V3�;�u>�E�Pj^VhH�V�X���t����E�PVhD�VW�\����J  jX��V��u�u�u�u�u�X��(  ���  9}u�V�EWWWW�u�uh   �u������u�;���   �}���$��7����e�ĉE�VWP�w������M���jXËe�3��}ԃM���u�9}���   WWV�u��u�uh   �u�������   �E�   �D6��$�������e�܉]��jXËe�3�3ۃM��;�tU�E;�u�V�M�<	�4f���f�N���S�u��u��uP�\��E�f�~���tf�>��uWS�u��/�����E��3��eȋM�d�    _^[��U��}
u�} }jj
�j �u�u�u�   �E��]�U��} �MSVWt�u�-A����u����3��u�Ƌ�3��u��	��v��W���0�A��wڀ! I����IG;�r�_^[]�������������U��WVS�u�}� V�x u;����
�t.�F�'G8�t�,A<ɀ� �A��,A<ɀ� �A8�t������x��`X�=\X j ���`Xj��S���$   ��   3ې
�t'�F�G8�t�PS�����؃�������8�t�������X�u	��`X�
j��S������[^_��U��WVS�M���   �u�}� V�x uN�A�Z� �I �&
�t!
�tFG8�r8�w�8�r8�w�8�uIu�3�8���   �������   ���   ��`X�=\X j ���`X��j��R���$   ��3�3ۋ����t#�tFGQPS�+����؃��!�����Y;�u	Iu�3�;�t	�����r��X�u	��`X���j��R�����ˋ�[^_��SUVW�|$�=P5~�jP����YY���\5�A����tG���7G��-��t��+u�7G3ۃ=P5~jV裬��YY��\5�p����t���\F��7G�σ�-��u��_^][�U��j�h��h�d�    Pd�%    ��SVW�e�TW3�;�u.WWjW�4���tj�WWjW�@�����   jX�TW��u�u�u�u�u�4��   ��u9}u�V�EWW�u�u�@��E�;�t]�}���$������e��u��jXËe�3�3��M��;�t3�u�V�u�u�@���t9}uWW��u�uj�Vj�u�̐�3��eЋM�d�    _^[��U��j�h�h�d�    Pd�%    ��SVW�e�XW3�;�u.VVjV�4���tj�VVjV�@�����   jX�XW��u�u�u�u�u�@��   ����   9uu�V�EVV�u�u�4��E�;�td�u����$������e���}��jXËe�3�3��M��;�t8�u�W�u�u�4���t$9uVVuVV��u�uj�Wh   �u����3��eЋM�d�    _^[����̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� V�t$��tV�}N��@P�1<��Y��YtVP�yM��YY^�3�^�̸T���  ��,�ES���A�I#�to3�8]tSS�2����Vt�T�����@�u�0��ES�M�E��)��V�N��YPV�M��v  �E�M�P�]��%   �E�h�P�E�$��1��^�M�[d�    �� �h��J  QQSV�E�W��P�u��E�I��,���]�e� �~j ��ψ����5����j S��!���M��h���_^[d�    �� �A��u����U���Q�M��g   �E�hX�P�1���|��  QV��u��h��e� j�N�1���M�����,���M�^d�    ��V�������D$tV�T��Y��^� ����c  QS�]VW��S�u��,���C�e� ���~j �ψ�����5����j S�� ���M��h���_^[d�    �� ����  QV��u��h��e� j�N�{���M������+���M�^d�    ��U���Q�M��*   �E�h�P�0��V�������D$tV���Y��^� V���t$�!����$���^� ����x
  QV��u��x��F$�e� ��v���W�F$���W ����   �N �����M�^d�    ��VW���w��t�vW�t$�V�6����_^� U��QV��M��$  �~$s�F$��dW��t;�t	@���F$r�F$�M��4�dW�v$���W�  ^��V��W3��N ;�t�&   WW�Ή~�F  �F   �~�~�~����_^�U��QV���Q  �M���   ��W�9���M��   ��^��VW��j �����F��t�8P�"����Y��u�F�f ��t�8P�����Y��u�f _^�j����VW�|$j��W�����tW�t$�v�Qh���F���~�$8 ��_^� ��WSVWj��_;�uh�W�Z����Wu5jh�W�P���uS��h���/��Y�=�W�%;�u�=�W�=�Wu
j�А��9=�WuS����_^[�jh�W�P���uh�W��Ã=�Wuh�W��øЍ�"  ��0�E�Vj �M��E�������V�sI��YPV�M�������e� �E�P�M��   �E�hX�P�EĀ��)-��^����  QQSV�E�W��P�u��E�I�?(���]�e� �~j ��ψ�'���5����j S�G���M������_^[d�    �� U���Q�M��g   �E�hȯP�,������G  QV��u�����e� j�N����M�����9(���M�^d�    ��V�������D$tV����Y��^� ����  QS�]VW��S�u��'���C�e� ���~j �ψ�T���5����j S�t���M������_^[d�    �� � ��  QV��u�����e� j�N����M�����'���M�^d�    ��U���Q�M��*   �E�hX�P�+��V�������D$tV���Y��^� V���t$�!��������^� �4��  ��0�E�Vj �M��E�������V�TG��YPV�M�������e� �E�P�M�������E�h��P�Eİ��
+��^�H��  QV��u�����e� j�N����M�����&���M�^d�    ��U���Q�M��*   �E�h��P�*��V�������D$tV�$��Y��^� V���t$�9��������^� �TXu�TX�   ��ku��k�   h@� �:,��Y�hm��.,��Y��2���   �   �h���,��Yù�W����U��QV��M��������M;Hs�P�4��3���u �} t�x t��W;Hs�@�4��3��M��.�����^�� U��QSV��M��{������W;�t2�8Xt
9�Wu��M��������^[�øf��#  QQV�M��;����e� �=�W ��   j(���Y�ȉM���E�t	j ��   �3��e� Wh���W�+����W��V�@?   ��W�x�$E��YYPV��������W��W�h����W_��t
��W��W�5�W�M���M��1����M��^d�    �øx��Y  Q�M��s�����W�e� ��t�]�����t�j����M���M�������M�d�    �ø���  QSV��W�u��F   ���M3��N�M�~�F�F�F�P�ωE��e���اS�:D��YPS�������M�����_^[d�    �� ���V���   �D$tV�k��Y��^� ����z  QQV��W�u����M��E�   �����~�E���v�FO����t��a�����t�j������v��+��Y�E��M�������e� j�N�
���M���_^d�    ���TXu�TX�   ��ku��k�   h@� �)��Y�hm��)��Yø��  QQ�ESV��3�WS�u��)
���E�NS�]���
���E�~ S���E���
���E�N0S�E����	��SS�E��ݿ��P�E��B������P�u��.���9]t�uS踿��Y;�Y��u�اW�B��YPW�N0�����M��_^[d�    �� ����   QV��u��F(�E�   ��v�F$��u���Pj �T���YYj�N0�R	��j�N �E��D	���e� j�N�6	���M��j���)	���M�^d�    ���TXu�TX�   ��ku��k�   h@� �'��Y�hm��'��Y���ku��k�    hm��t'��Y��TXu�TX�    h@� �S'��Y��%ܐ��j�Pd�    P�D$d�%    �l$�l$P�̋D$��tD�T$VW��|$׃�t2�   t�:uRFGHt��8�uE�N�W8�u;������u�_^Ëȃ���t+�t'�N��W�8�u8�u����8�u8��    �_���^Å�tċ�8�u�Ht8�u�Ht��  � ��  � ;�u�H_^����̸���7!�������̸��'!�������̸@��!���̍M����������!���̋M��  ��� ��� ���̋M������h��� ���̋M���������� ���̋M��������� ���̋M��� �������� ����̍M��f����h�� ���̋M��������s ���̋M��p���د�_ ���̋M��\��� ��K ���̋M��H���(��7 ���̍M���������# ���̋M�� ������ ���̍M������u�����Yø������M������������̋M������8������̋M��	����M�������M��\����`������̋M��n����M���c����M�� �X����M��0�M�������n��̋M��:����M����/����M��� �$����ر�E��                                                                                                                                                                                                                                    8� $� T�     �� |�     �� �� ʵ     �  � "� � �� � Ҽ ¼ �� �� �� �� n� ޴ H� <� 2� &� � � �� � һ » �� �� �� l� T� >� $� 
� �� � ں Ⱥ �� �� δ �� X� �� �� �� �� �� �� �� ĸ и ޸ � � � &� 8� L� h� �� �� �� ƹ Թ � � �� � &� 2� >� T� n� ~� 4�     � � �� � ܷ ̷ �� �� �� �� �� z� j� V� F� 6� &� � �� � Զ ƶ �� �� �� �� ~� t� d� R� F� 4�  � � ��     ^� J� 8� 0�  �     t�             H�z��o@      �?      �?     �o@               @-�-n0_�?q���h �?      �?      Y@���(\�_�UUUUU�?���m0_�?���m0_�?    �< �; ������@= �= �= A ���> p��A pA ��pB �H �� C Љ�G �H P�0�`�D p�pG p� �0�����@�P�P��B P�P�P��< ����P�ЉP� �P�0�`�`�p� �p� �0�����@�P�P�P�P�P�P��.eB0Q }�}�}�}�}� R pZ �l �[  e P� � `� �� �� Ћ �� ��  � �� `� �� �� Ћ �    Г P� �� �� Ћ  � ��  � �� p� � �� Ћ �0�     P       �h㈵��>      �?�e Pi �i j Pj `� �l �l P� �l �k P��l �l �l Pp �l �p P��l �l �l q �q �r s �l �l �l Ps �l  t P��l pt �l P� �l @z pz �l   �?�l �l �{ �q �}  � �l �l �l  ~ �q �  � @� �l �l P� �l �� P��l Ђ �l @� �q @� P��l �l �l �l p� �q Ѕ  � �l ����       �� �� �� 0� �< ����P�ЉP� �P�0�`�`�p� � p�p�����p� �����Љ����p����l Ўp������P�P���    ����MbP?�������?      �?     �r@      y@�}�P�p!�!P(������0,�(0�Љ��Ќ -�-��Љ��Љp���`-��}��.�-��Љ��Љp���`-���.�0�-�0Љ��Љp��1`-���00�����Љ��Љp����l �� �������P���0�Љ��Ќ������Љ��Љp����l Ў   O  zD�< �� �p�����P�P���p�Ŭ~�Unknown exception   ����csm�               �        ����    ]�����    ������    _�����    ������     �����    |�   �~PA   ���GAIsProcessorFeaturePresent   KERNEL32    e+000         �?5�h!���>@�������             ��      �@      �            ��������    ����    �    �������U�Y�    ��������    ����    $�    ������    z�    f�j�       EEE50 P     (8PX 700WP        `h````  ppxxxx          ( n u l l )     (null)      ����    l�����    ��__GLOBAL_HEAP_SELECTED  __MSVCRT_HEAP_SELECT    runtime error   
  TLOSS error
   SING error
    DOMAIN error
  R6028
- unable to initialize heap
    R6027
- not enough space for lowio initialization
    R6026
- not enough space for stdio initialization
    R6025
- pure virtual function call
   R6024
- not enough space for _onexit/atexit table
    R6019
- unable to open console device
    R6018
- unexpected heap error
    R6017
- unexpected multithread lock error
    R6016
- not enough space for thread data
 
abnormal program termination
    R6009
- not enough space for environment
 R6008
- not enough space for arguments
   R6002
- floating point not loaded
    Microsoft Visual C++ Runtime Library    

  Runtime Error!

Program:    <program name unknown>  _yn _y1 _y0 frexp   fmod    _hypot  _cabs   ldexp   modf    fabs    floor   ceil    tan cos sin sqrt    atan2   atan    acos    asin    tanh    cosh    sinh    log10   log pow exp �������             ��      �@      �        ����    3����    �3GetLastActivePopup  GetActiveWindow MessageBoxA user32.dll              �����J�JLC_TIME LC_NUMERIC  LC_MONETARY LC_CTYPE    LC_COLLATE  LC_ALL  ;   =;  =   _., .   _       ����\R`R����SS1#QNAN  1#INF   1#IND   1#SNAN  Paraguay    Uruguay Chile   Ecuador Argentina   Peru    Colombia    Venezuela   Dominican Republic  South Africa    Panama  Luxembourg  Costa Rica  Switzerland Guatemala   Canada  Spanish - Modern Sort   Australia   English Austria German  Belgium Mexico  Spanish Basque  Sweden  Swedish Iceland Icelandic   France  French  Finland Finnish Spain   Spanish - Traditional Sort  united-states   united-kingdom  trinidad & tobago   south-korea south-africa    south korea south africa    slovak  puerto-rico pr-china    pr china    nz  new-zealand hong-kong   holland great britain   england czech   china   britain america usa us  uk  swiss   swedish-finland spanish-venezuela   spanish-uruguay spanish-puerto rico spanish-peru    spanish-paraguay    spanish-panama  spanish-nicaragua   spanish-modern  spanish-mexican spanish-honduras    spanish-guatemala   spanish-el salvador spanish-ecuador spanish-dominican republic  spanish-costa rica  spanish-colombia    spanish-chile   spanish-bolivia spanish-argentina   portuguese-brazilian    norwegian-nynorsk   norwegian-bokmal    norwegian   italian-swiss   irish-english   german-swiss    german-luxembourg   german-lichtenstein german-austrian french-swiss    french-luxembourg   french-canadian french-belgian  english-usa english-us  english-uk  english-trinidad y tobago   english-south africa    english-nz  english-jamaica english-ire english-caribbean   english-can english-belize  english-aus english-american    dutch-belgian   chinese-traditional chinese-singapore   chinese-simplified  chinese-hongkong    chinese chi chh canadian    belgian australian  american-english    american english    american    OCP ACP H:mm:ss dddd, MMMM dd, yyyy M/d/yy  PM  AM  December    November    October September   August  July    June    April   March   February    January Dec Nov Oct Sep Aug Jul Jun May Apr Mar Feb Jan Saturday    Friday  Thursday    Wednesday   Tuesday Monday  Sunday  Sat Fri Thu Wed Tue Mon Sun     ����yy����_ycySunMonTueWedThuFriSat   JanFebMarAprMayJunJulAugSepOctNovDec    �����}�}    �����~�~             ���`�}�ios::eofbit set ios::failbit set    ios::badbit set X�ǀ`�m����p ��`��string too long @�<�`������`�چinvalid string position    *   (������� ȫ�� 0� @� P�  � � x��� � � @� P� `� � ��� ~�p�         ��        ����        @�               X�            ��`�            ����        ��               ��            ��    H       ����        0H       ����        �Ш@�                �            0H�    Ш@�                   8�            HH�    XH        ����        p�               ��            XH��    xH       ����        �H       ����        Щ��@�               �            �H��    ��@�                    �            xH0�    �H       ����        X���@�               p�            �H��ت                   ��            �H��    �H        ����        �H       ����        �ت                   �            �H�     I       ����        @�ت                   X�             Ih�    xI       ����        ��ت                   ��            xI��    ��       ����        �@�                   ��            ���        ��    ����       �        ��    ����       Њ        P�0�        `�     p� �   ��   ��            ����    ����                  ج                m�  �   �   �            ����    ����                  0�                ��  �   `�   p�            ����    ����                  ��                �     H    ����       �        0H    ����       ��       ����0�    @�    ح �   �                    ����L� �   @�                    ����`�   ��0�        ��    H� �   ��                    ����t� �   ��                    ������ �   خ                    ������ �    �                    ������    xH    ����       X�        �H    ����       +�       (��0�    ��    H� �   ��                    ����ȍ �   ��                    ����܍   �0�        ��    �� �   ��                    ������ �    �                    ����� �   H�                    �����    �H    ����       �       P��0�    ��    p� �   ��                    ����,� �   ذ                    ����@� �    �                    ����T�    \� �   0�                    ����p� �   X�                    ������ �   ��                    ������    ��   �� �   ��                    ������    Ȏ   ӎ   ގ �   ��                    �����    ��   �ܲ         � ,� ��         p� � ��         �� � ̲         ޵ � �         � X� ��         d�  � ��         ��  �                     8� $� T�     �� |�     �� �� ʵ     �  � "� � �� � Ҽ ¼ �� �� �� �� n� ޴ H� <� 2� &� � � �� � һ » �� �� �� l� T� >� $� 
� �� � ں Ⱥ �� �� δ �� X� �� �� �� �� �� �� �� ĸ и ޸ � � � &� 8� L� h� �� �� �� ƹ Թ � � �� � &� 2� >� T� n� ~� 4�     � � �� � ܷ ̷ �� �� �� �� �� z� j� V� F� 6� &� � �� � Զ ƶ �� �� �� �� ~� t� d� R� F� 4�  � � ��     ^� J� 8� 0�  �     t�     �Sleep  CloseHandle J CreateThread  � FormatMessageA  GetLastError  D CreateProcessA  KERNEL32.dll  � DestroyWindow � GetDC Y CreateWindowExA �RegisterClassExA  � DefWindowProcA  USER32.dll  �SetPixelFormat   ChoosePixelFormat GDI32.dll  gluLookAt   gluPerspective   gluBuild2DMipmaps GLU32.dll ZwglCreateContext  j glGenTextures C glDeleteTextures  \wglDeleteContext  ewglMakeCurrent  glScaled  � glLoadIdentity  � glMatrixMode   glClear WglViewport  P glEnable  a glFinish  8glTexParameteri  glBindTexture � glPopMatrix H glDisableClientState  K glDrawElements  VglVertexPointer Q glEnableClientState � glMultMatrixf � glPushMatrix  4glTexImage1D  dwglGetProcAddress 5glTexImage2D  )glTexCoordPointer � glNormalPointer R glEnd >glVertex2d   glBegin * glColor4d  glClearColor  � glHint  � glReadPixels  `wglGetCurrentDC } glGetString OPENGL32.dll   CgFXCreateEffect   CgFXCreateEffectFromFileA  CgFXSetDevice CgFXParser.dll  � timeGetTime WINMM.dll /RtlUnwind RaiseException  �HeapFree  �HeapReAlloc �HeapAlloc } ExitProcess �TerminateProcess  � GetCurrentProcess � GetCommandLineA tGetVersion  >GetProcAddress  &GetModuleHandleA  �InitializeCriticalSection U DeleteCriticalSection f EnterCriticalSection  �LeaveCriticalSection  � GetCurrentThreadId  �TlsSetValue �TlsAlloc  �TlsFree qSetLastError  �TlsGetValue �SetUnhandledExceptionFilter �HeapSize  ReadFile  $GetModuleFileNameA  	GetEnvironmentVariableA uGetVersionExA �HeapDestroy �HeapCreate  �VirtualFree �VirtualAlloc  �IsBadWritePtr mSetHandleCount  RGetStdHandle  GetFileType PGetStartupInfoA � FreeEnvironmentStringsA � FreeEnvironmentStringsW �WideCharToMultiByte GetEnvironmentStrings GetEnvironmentStringsW  �WriteFile �InterlockedDecrement  �InterlockedIncrement  �IsBadReadPtr  �IsBadCodePtr  jSetFilePointer  |SetStdHandle  � FlushFileBuffers  4 CreateFileA � GetCPInfo � GetACP  1GetOEMCP  �LoadLibraryA  �MultiByteToWideChar SGetStringTypeA  VGetStringTypeW  �LCMapStringA  �LCMapStringW  aSetEndOfFile  �IsValidLocale �IsValidCodePage GetLocaleInfoA  w EnumSystemLocalesA  qGetUserDefaultLCID  GetLocaleInfoW  �InterlockedExchange           !@    ��          x� |� �� �� ��   c4dfx.cdl c4d_main                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �� @
����+�q�T�ċ�'�        ����'F��        ��        ��    C:\Dokumente und Einstellungen\jl.2G5\Desktop\C4D 8.5, SketchAndToon\8500\030911 8.500\plugins\c4dfx\source\BitmapWrapper.cpp   C4Dfx:      C:\Dokumente und Einstellungen\jl.2G5\Desktop\C4D 8.5, SketchAndToon\8500\030911 8.500\plugins\c4dfx\source\C4DWrapper.cpp  Camera is not in perspective mode.  C:\Dokumente und Einstellungen\jl.2G5\Desktop\C4D 8.5, SketchAndToon\8500\030911 8.500\plugins\c4dfx\source\FXCommand.cpp   fx32.tif    ... Could not open window.  Could not allocate window.  C:\Dokumente und Einstellungen\jl.2G5\Desktop\C4D 8.5, SketchAndToon\8500\030911 8.500\plugins\c4dfx\source\FXDialog.cpp    C:\Dokumente und Einstellungen\jl.2G5\Desktop\C4D 8.5, SketchAndToon\8500\030911 8.500\plugins\c4dfx\source\FXMaterial.cpp  Edit .fx file?  Mfxmaterial Shadows: No suitable OpenGL format found.   Shadows: Coudn't create render context. Shadows: Couldn't create device context.    Shadows: Couldn't create depth buffer.  Isn't a polygon object (in computation of shadow map).  );
	}
} ,
			lightPos   , lightCol  , lightParams   , lightUp   , lightDir  , lightSide 			lumiCol, diffCol, bumpHeight, enviCol, specCol   			depthSampler 	OUT.col = colorSum;
	return OUT;
}
technique t0
{
	pass p0
	{
		VertexShader = compile vs_2_x mainVS(wvp, wit, w, vit);
		ZEnable = true;
		ZWriteEnable = true;
		CullMode = None;
		PixelShader = compile ps_2_x mainPS(diffuseSampler, specShapeSampler, normalSampler, envMapSampler,
 		colorSum += shadowFactor*baseCol*lightCol .rgb;
	}
   		float d = dot(Ld, lightDir    .xyz);
		float z = 10.1010101/d + 1.01010101;
		float2 depthUV = float2(0.5, 0.5) + 0.5*float2(dot(L1, lightSide    .xyz), dot(L1, lightUp  .xyz));
		shadowFactor *= max(lightParams   .y, tex2Dproj(depthSampler  , float4(depthUV.x, depthUV.y, z-0.0002, 1.0)).x);
 	{
		float3 Ld = lightPos   .xyz - IN.wPos;
		float3 Ln = normalize(Ld);
		float3 baseCol = max(0.0, dot(Ln, Nb))*baseDiffCol;
		float spec = tex1D(specShapeSampler, dot(Vn, reflect(Ln, Nb))).r;
		baseCol += specCol.rgb*spec;
		float3 L1 = (Ln/dot(Ln, lightDir    .xyz) - lightDir    .xyz)*lightParams   .z;
		float shadowFactor = max(lightParams  .x, smoothstep(1.0, lightParams .w, length(L1)));
  )
{
	pixelOutput OUT;
	float3 Vn = normalize(IN.view);
	float3 Nn = normalize(IN.norm);
	float3 tangn = normalize(IN.tang);
	float3 binormn = normalize(IN.binorm);
	float2 bumps = bumpHeight*(tex2D(normalSampler, IN.uv.xy).xy * 2.0 - float2(1.0, 1.0));
	float3 Nb = normalize(bumps.x*tangn + bumps.y*binormn + Nn);
	float3 env = texCUBE(enviSampler, reflect(Vn, Nb)).rgb;
	float3 colorSum = lumiCol.rgb + env*enviCol.rgb;
	float3 baseDiffCol = diffCol.rgb + tex2D(diffuseSampler, IN.uv.xy).rgb;
 ,
	uniform float4 lightPos  ,
	uniform float4 lightCol  ,
	uniform float4 lightParams   ,
	uniform float4 lightUp   ,
	uniform float4 lightDir  ,
	uniform float4 lightSide 	uniform float4 lumiCol,
	uniform float4 diffCol,
	uniform float bumpHeight,
	uniform float4 enviCol,
	uniform float4 specCol   	uniform sampler2D depthSampler ,
  struct appdata {
	float4 position	: POSITION;
	float4 norm : NORMAL;
	float4 uv: TEXCOORD0;
	float4 tang : TEXCOORD1;
	float4 binorm : TEXCOORD2;
};
struct vertexOutput {
	float4 hPos : POSITION;
	float4 uv : TEXCOORD0;
	float3 norm : TEXCOORD1;
	float3 tang : TEXCOORD2;
	float3 binorm : TEXCOORD3;
	float3 view : TEXCOORD4;
	float3 wPos : TEXCOORD5;
};
struct pixelOutput {
	float3 col : COLOR;
};
vertexOutput mainVS(appdata IN,
	uniform float4x4 wvp,
	uniform float4x4 wit,
	uniform float4x4 w,
	uniform float4x4 vit)
{
	vertexOutput OUT;
	OUT.uv = IN.uv;
	OUT.hPos = mul(wvp, IN.position);
	OUT.norm = mul(wit, IN.norm).xyz;
	OUT.tang = mul(w, IN.tang).xyz;
	OUT.binorm = mul(w, IN.binorm).xyz;
	float3 pW = mul(w, IN.position).xyz;
	OUT.wPos = pW;
	OUT.view = normalize(pW - vit[3].xyz);
	return OUT;
}
pixelOutput mainPS(vertexOutput IN,
	uniform sampler2D diffuseSampler,
	uniform sampler1D specShapeSampler,
	uniform sampler2D normalSampler,
	uniform samplerCUBE enviSampler,
   sampler2D depthSampler   = sampler_state
{	Texture = <depthTexture  >;
	MinFilter = Linear;
	MagFilter = Linear;
	MipFilter = None;
	AddressU = Border;
	AddressV = Border;
	BorderColor = {0.0f, 0.0f, 0.0f, 1.0f};
};
    sampler2D diffuseSampler = sampler_state
{	Texture = <diffuseTexture>;
	MinFilter = Linear;
	MagFilter = Linear;
	MipFilter = Linear;
};
sampler1D specShapeSampler = sampler_state
{	Texture = <specShapeTexture>;
	AddressU = Clamp;
	MinFilter = Linear;
	MagFilter = Linear;
	MipFilter = None;
};
sampler2D normalSampler = sampler_state
{	Texture = <normalTexture>;
	MinFilter = Linear;
	MagFilter = Linear;
	MipFilter = Linear;
};
samplerCUBE envMapSampler = sampler_state
{	Texture = <enviTexture>;
	MinFilter = Linear;
	MagFilter = Linear;
	MipFilter = Linear;
};
   texture depthTexture    float4 lightPos ;
float4 lightCol   ;
float4 lightParams    ;
float4 lightUp    ;
float4 lightDir   ;
float4 lightSide  ;
  float4x4 wvp;
float4x4 wit;
float4x4 w;
float4x4 vit;
float4 diffCol;
float4 lumiCol;
texture diffuseTexture;
float bumpHeight;
texture normalTexture;
float4 enviCol;
texture enviTexture;
texture specShapeTexture;
float4 specCol;
  --- Object  Desc    Couldn't allocate parameter.    UNKNOWN TYPE    slider  gui uistep  uimax   uimin   WorldViewProjectionIT   WorldViewProjectionT    WorldViewProjectionI    WorldViewProjection ProjectionIT    ProjectionT ProjectionI Projection  WorldViewIT WorldViewT  WorldViewI  WorldView   ViewIT  ViewT   ViewI   View    WorldIT WorldT  WorldI  World   Emissive    Specular    Diffuse Ambient default File    Couldn't load:  No .dds file:   .dds    No object linked for position or direction parameter?   Space   DIRECTION   POSITION        ��    .?AVexception@@ ��    .?AVbad_cast@std@@  missing locale facet    C   ,   e   E   %p  true    false   Shadows: Allocation error.  C:\Dokumente und Einstellungen\jl.2G5\Desktop\C4D 8.5, SketchAndToon\8500\030911 8.500\plugins\c4dfx\source\LightsMaterialsObjects.cpp  Materials: Allocation error.    error on reading    error on setting and validating technique   error on retrieving FXWrapper   error on retrieving technique   error on setting and validating emulator technique  error on loading emulator fx    C4Dfx: material     No standard or C4Dfx material.  Couldn't retrieve Cast Shadow setting   Tlight  fx24.tif    C:\Dokumente und Einstellungen\jl.2G5\Desktop\C4D 8.5, SketchAndToon\8500\030911 8.500\plugins\c4dfx\source\LightTag.cpp    This version of C4Dfx needs Cinema 4D 8.5 or later. DDS     rb  glCompressedTexImage1DARB   glCompressedTexImage2DARB   glTexImage3D    glCompressedTexImage3DARB   Couldn't allocate memory.   CgFX: pass failed.  Effect initialization failed.   uvw tag inaccessible.   Isn't a polygon object. No standard material or faulty C4Dfx material.  C:\Dokumente und Einstellungen\jl.2G5\Desktop\C4D 8.5, SketchAndToon\8500\030911 8.500\plugins\c4dfx\source\PrefDialog.cpp  /L:<LINE> "<FILE>"  C4Dfx.prefs <FILE>  <LINE>  %8.3f s No suitable OpenGL format found.    Couldn't allocate materials.    Couldn't allocate shadows.  Couldn't allocate lights.   Switching CgFX to OpenGL device failed. OpenGL  Couldn't switch to offscreen render context.    Couldn't create offscreen render context.   Couldn't create device context. Couldn't create offscreen buffer.   Couldn't open movie file.   Couldn't allocate output bitmap.    No path specified for saving output.    Only user-defined AVI can be used as output format. Couldn't allocate memory for double buffering.  Couldn't allocate memory for renderer.  Couldn't write frame to movie.  Couldn't switch back to main render context.    Could not create renderer thread.   Could not initialize renderer context.  Could not allocate renderer.    Could not create renderer window.   C4Dfx   Failing due to error on program startup.    Couldn't switch back to offscreen render context.   C4dfx:   frames finished    C4dfx: frame     of     Rendering ...   Couldn't attach preview area.   Couldn't create preview area.   Couldn't open preview window.   Couldn't start rendering thread.    Couldn't create rendering thread.   C:\Dokumente und Einstellungen\jl.2G5\Desktop\C4D 8.5, SketchAndToon\8500\030911 8.500\plugins\c4dfx\source\RenderDialog.cpp    Couldn't clone document for rendering.  Couldn't open renderer window.  (  $                                   GL_NV_multisample_filter_hint   Driver does not support WGL_NV_render_depth_texture WGL_ARB_render_texture  GL_ARB_depth_texture    WGL_ARB_pbuffer WGL_ARB_pixel_format    GL_ARB_multisample  GL_ARB_multitexture WGL_ARB_extensions_string   Not support of wglGetProcAddress. Use vendor specific driver?   Couldn't switch to rendering context for initial window.    Couldn't create rendering context for initial window.   Couldn't set OpenGL pixel format for initial window.    No suitable OpenGL pixel format for initial window. Couldn't get device context of initial window.  Couldn't create initial window. Couldn't register window class. Cannot open editor:
    WGL_NV_render_texture_rectangle WGL_NV_float_buffer wglGetSwapIntervalEXT   wglSwapIntervalEXT  WGL_EXT_swap_control    wglGetExtensionsStringEXT   WGL_EXT_extensions_string   wglSetPbufferAttribARB  wglReleaseTexImageARB   wglBindTexImageARB  wglChoosePixelFormatARB wglGetPixelFormatAttribfvARB    wglGetPixelFormatAttribivARB    wglQueryPbufferARB  wglDestroyPbufferARB    wglReleasePbufferDCARB  wglGetPbufferDCARB  wglCreatePbufferARB wglGetExtensionsStringARB   wglRestoreBufferRegionARB   wglSaveBufferRegionARB  wglDeleteBufferRegionARB    wglCreateBufferRegionARB    WGL_ARB_buffer_region   GL_SGIX_shadow  GL_SGIX_depth_texture   GL_SGIS_texture_lod GL_SGIS_generate_mipmap GL_NV_vertex_program2   GL_NV_vertex_program1_1 glVertexAttribs4ubvNV   glVertexAttribs4svNV    glVertexAttribs4fvNV    glVertexAttribs4dvNV    glVertexAttribs3svNV    glVertexAttribs3fvNV    glVertexAttribs3dvNV    glVertexAttribs2svNV    glVertexAttribs2fvNV    glVertexAttribs2dvNV    glVertexAttribs1svNV    glVertexAttribs1fvNV    glVertexAttribs1dvNV    glVertexAttrib4ubvNV    glVertexAttrib4svNV glVertexAttrib4sNV  glVertexAttrib4fvNV glVertexAttrib4fNV  glVertexAttrib4dvNV glVertexAttrib4dNV  glVertexAttrib3svNV glVertexAttrib3sNV  glVertexAttrib3fvNV glVertexAttrib3fNV  glVertexAttrib3dvNV glVertexAttrib3dNV  glVertexAttrib2svNV glVertexAttrib2sNV  glVertexAttrib2fvNV glVertexAttrib2fNV  glVertexAttrib2dvNV glVertexAttrib2dNV  glVertexAttrib1svNV glVertexAttrib1sNV  glVertexAttrib1fvNV glVertexAttrib1fNV  glVertexAttrib1dvNV glVertexAttrib1dNV  glVertexAttribPointerNV glTrackMatrixNV glRequestResidentProgramsNV glProgramParameters4fvNV    glProgramParameters4dvNV    glProgramParameter4fvNV glProgramParameter4fNV  glProgramParameter4dvNV glProgramParameter4dNV  glLoadProgramNV glIsProgramNV   glGetVertexAttribPointervNV glGetVertexAttribivNV   glGetVertexAttribfvNV   glGetVertexAttribdvNV   glGetTrackMatrixivNV    glGetProgramStringNV    glGetProgramivNV    glGetProgramParameterfvNV   glGetProgramParameterdvNV   glGenProgramsNV glExecuteProgramNV  glDeleteProgramsNV  glBindProgramNV glAreProgramsResidentNV GL_NV_vertex_program    GL_NV_vertex_array_range2   wglFreeMemoryNV wglAllocateMemoryNV glVertexArrayRangeNV    glFlushVertexArrayRangeNV   GL_NV_vertex_array_range    GL_NV_texture_shader3   GL_NV_texture_shader2   GL_NV_texture_shader    GL_NV_texture_rectangle GL_NV_texture_env_combine4  GL_NV_texture_compression_vtc   GL_NV_texgen_reflection glActiveStencilFaceNV   GL_NV_stencil_two_side  glGetCombinerStageParameterfvNV glCombinerStageParameterfvNV    GL_NV_register_combiners2   glGetFinalCombinerInputParameterivNV    glGetFinalCombinerInputParameterfvNV    glGetCombinerOutputParameterivNV    glGetCombinerOutputParameterfvNV    glGetCombinerInputParameterivNV glGetCombinerInputParameterfvNV glFinalCombinerInputNV  glCombinerOutputNV  glCombinerInputNV   glCombinerParameteriNV  glCombinerParameterivNV glCombinerParameterfNV  glCombinerParameterfvNV GL_NV_register_combiners    glPrimitiveRestartIndexNV   glPrimitiveRestartNV    GL_NV_primitive_restart glPointParameterivNV    glPointParameteriNV GL_NV_point_sprite  glFlushPixelDataRangeNV glPixelDataRangeNV  GL_NV_pixel_data_range  GL_NV_packed_depth_stencil  glGetOcclusionQueryuivNV    glGetOcclusionQueryivNV glEndOcclusionQueryNV   glBeginOcclusionQueryNV glIsOcclusionQueryNV    glDeleteOcclusionQueriesNV  glGenOcclusionQueriesNV GL_NV_occlusion_query   GL_NV_light_max_exponent    glVertexAttribs4hvNV    glVertexAttribs3hvNV    glVertexAttribs2hvNV    glVertexAttribs1hvNV    glVertexAttrib4hvNV glVertexAttrib4hNV  glVertexAttrib3hvNV glVertexAttrib3hNV  glVertexAttrib2hvNV glVertexAttrib2hNV  glVertexAttrib1hvNV glVertexAttrib1hNV  glVertexWeighthvNV  glVertexWeighthNV   glSecondaryColor3hvNV   glSecondaryColor3hNV    glFogCoordhvNV  glFogCoordhNV   glMultiTexCoord4hvNV    glMultiTexCoord4hNV glMultiTexCoord3hvNV    glMultiTexCoord3hNV glMultiTexCoord2hvNV    glMultiTexCoord2hNV glMultiTexCoord1hvNV    glMultiTexCoord1hNV glTexCoord4hvNV glTexCoord4hNV  glTexCoord3hvNV glTexCoord3hNV  glTexCoord2hvNV glTexCoord2hNV  glTexCoord1hvNV glTexCoord1hNV  glColor4hvNV    glColor4hNV glColor3hvNV    glColor3hNV glNormal3hvNV   glNormal3hNV    glVertex4hvNV   glVertex4hNV    glVertex3hvNV   glVertex3hNV    glVertex2hvNV   glVertex2hNV    GL_NV_half_float    glGetProgramNamedParameterdvNV  glGetProgramNamedParameterfvNV  glProgramNamedParameter4dvNV    glProgramNamedParameter4fvNV    glProgramNamedParameter4dNV glProgramNamedParameter4fNV GL_NV_fragment_program  GL_NV_fog_distance  GL_NV_float_buffer  glGetFenceivNV  glIsFenceNV glFinishFenceNV glTestFenceNV   glSetFenceNV    glDeleteFencesNV    glGenFencesNV   GL_NV_fence glMultiDrawRangeElementArrayNV  glMultiDrawElementArrayNV   glDrawRangeElementArrayNV   glDrawElementArrayNV    glElementPointerNV  GL_NV_element_array GL_NV_depth_clamp   GL_NV_copy_depth_to_color   GL_NV_blend_square  GL_IBM_texture_mirrored_repeat  GL_HP_occlusion_test    glVertexWeightPointerEXT    glVertexWeightfvEXT glVertexWeightfEXT  GL_EXT_vertex_weighting glDrawArraysEXT glVertexPointerEXT  glTexCoordPointerEXT    glNormalPointerEXT  glIndexPointerEXT   glGetPointervEXT    glEdgeFlagPointerEXT    glColorPointerEXT   glArrayElementEXT   GL_EXT_vertex_array glTexImage3DEXT GL_EXT_texture3D    glPrioritizeTexturesEXT glIsTextureEXT  glGenTexturesEXT    glDeleteTexturesEXT glBindTextureEXT    glAreTexturesResidentEXT    GL_EXT_texture_object   GL_EXT_texture_lod_bias GL_EXT_texture_filter_anisotropic   GL_EXT_texture_env_dot3 GL_EXT_texture_env_combine  GL_EXT_texture_env_add  GL_EXT_texture_compression_s3tc GL_EXT_stencil_wrap glActiveStencilFaceEXT  GL_EXT_stencil_two_side GL_EXT_shared_texture_palette   GL_EXT_shadow_funcs GL_EXT_separate_specular_color  glSecondaryColorPointerEXT  glSecondaryColor3usvEXT glSecondaryColor3usEXT  glSecondaryColor3uivEXT glSecondaryColor3uiEXT  glSecondaryColor3ubvEXT glSecondaryColor3ubEXT  glSecondaryColor3svEXT  glSecondaryColor3sEXT   glSecondaryColor3ivEXT  glSecondaryColor3iEXT   glSecondaryColor3fvEXT  glSecondaryColor3fEXT   glSecondaryColor3dvEXT  glSecondaryColor3dEXT   glSecondaryColor3bvEXT  glSecondaryColor3bEXT   GL_EXT_secondary_color  GL_EXT_rescale_normal   glPointParameterfvEXT   glPointParameterfEXT    GL_EXT_point_parameters glGetColorTableParameterivEXT   glGetColorTableParameterfvEXT   glGetColorTableEXT  glColorTableEXT glColorSubTableEXT  GL_EXT_paletted_texture GL_EXT_packed_pixels    glMultiDrawElementsEXT  glMultiDrawArraysEXT    GL_EXT_multi_draw_arrays    glFogCoordPointerEXT    glFogCoordfvEXT glFogCoordfEXT  glFogCoorddvEXT glFogCoorddEXT  GL_EXT_fog_coord    GL_EXT_draw_range_elements  glUnlockArraysEXT   glLockArraysEXT GL_EXT_compiled_vertex_array    GL_EXT_blend_subtract   glBlendEquationEXT  GL_EXT_blend_minmax glBlendFuncSeparateEXT  GL_EXT_blend_func_separate  glBlendColorEXT GL_EXT_blend_color  GL_EXT_bgra GL_EXT_abgr glWindowPos3svARB   glWindowPos3ivARB   glWindowPos3fvARB   glWindowPos3dvARB   glWindowPos3sARB    glWindowPos3iARB    glWindowPos3fARB    glWindowPos3dARB    glWindowPos2svARB   glWindowPos2ivARB   glWindowPos2fvARB   glWindowPos2dvARB   glWindowPos2sARB    glWindowPos2iARB    glWindowPos2fARB    glWindowPos2dARB    GL_ARB_window_pos   glIsProgramARB  glGetVertexAttribPointervARB    glGetVertexAttribivARB  glGetVertexAttribfvARB  glGetVertexAttribdvARB  glGetProgramStringARB   glGetProgramivARB   glGetProgramLocalParameterfvARB glGetProgramLocalParameterdvARB glGetProgramEnvParameterfvARB   glGetProgramEnvParameterdvARB   glProgramLocalParameter4fvARB   glProgramLocalParameter4fARB    glProgramLocalParameter4dvARB   glProgramLocalParameter4dARB    glProgramEnvParameter4fvARB glProgramEnvParameter4fARB  glProgramEnvParameter4dvARB glProgramEnvParameter4dARB  glGenProgramsARB    glDeleteProgramsARB glBindProgramARB    glProgramStringARB  glDisableVertexAttribArrayARB   glEnableVertexAttribArrayARB    glVertexAttribPointerARB    glVertexAttrib4NuivARB  glVertexAttrib4NusvARB  glVertexAttrib4NubvARB  glVertexAttrib4NivARB   glVertexAttrib4NsvARB   glVertexAttrib4NbvARB   glVertexAttrib4dvARB    glVertexAttrib4fvARB    glVertexAttrib4uivARB   glVertexAttrib4usvARB   glVertexAttrib4ubvARB   glVertexAttrib4ivARB    glVertexAttrib4svARB    glVertexAttrib4bvARB    glVertexAttrib3dvARB    glVertexAttrib3fvARB    glVertexAttrib3svARB    glVertexAttrib2dvARB    glVertexAttrib2fvARB    glVertexAttrib2svARB    glVertexAttrib1dvARB    glVertexAttrib1fvARB    glVertexAttrib1svARB    glVertexAttrib4NubARB   glVertexAttrib4dARB glVertexAttrib4fARB glVertexAttrib4sARB glVertexAttrib3dARB glVertexAttrib3fARB glVertexAttrib3sARB glVertexAttrib2dARB glVertexAttrib2fARB glVertexAttrib2sARB glVertexAttrib1dARB glVertexAttrib1fARB glVertexAttrib1sARB GL_ARB_vertex_program   glMultTransposeMatrixdARB   glMultTransposeMatrixfARB   glLoadTransposeMatrixdARB   glLoadTransposeMatrixfARB   GL_ARB_transpose_matrix GL_ARB_texture_mirrored_repeat  GL_ARB_texture_env_dot3 GL_ARB_texture_env_combine  GL_ARB_texture_env_add  GL_ARB_texture_cube_map glGetCompressedTexImageARB  glCompressedTexSubImage1DARB    glCompressedTexSubImage2DARB    glCompressedTexSubImage3DARB    GL_ARB_texture_compression  GL_ARB_texture_border_clamp GL_ARB_shadow   glPointParameterfvARB   glPointParameterfARB    GL_ARB_point_parameters glClientActiveTextureARB    glActiveTextureARB  glMultiTexCoord4svARB   glMultiTexCoord4sARB    glMultiTexCoord4ivARB   glMultiTexCoord4iARB    glMultiTexCoord4fvARB   glMultiTexCoord4fARB    glMultiTexCoord4dvARB   glMultiTexCoord4dARB    glMultiTexCoord3svARB   glMultiTexCoord3sARB    glMultiTexCoord3ivARB   glMultiTexCoord3iARB    glMultiTexCoord3fvARB   glMultiTexCoord3fARB    glMultiTexCoord3dvARB   glMultiTexCoord3dARB    glMultiTexCoord2svARB   glMultiTexCoord2sARB    glMultiTexCoord2ivARB   glMultiTexCoord2iARB    glMultiTexCoord2fvARB   glMultiTexCoord2fARB    glMultiTexCoord2dvARB   glMultiTexCoord2dARB    glMultiTexCoord1svARB   glMultiTexCoord1sARB    glMultiTexCoord1ivARB   glMultiTexCoord1iARB    glMultiTexCoord1fvARB   glMultiTexCoord1fARB    glMultiTexCoord1dvARB   glMultiTexCoord1dARB    GL_ARB_fragment_program Error allocating memory in file %s, line %d
    C:\Programme\Microsoft Visual Studio\VC98\INCLUDE\glh/glh_extensions.h  1.3 GL_VERSION_1_4  1.2 GL_VERSION_1_3  1.1 1.0 GL_VERSION_1_2  res C:\Dokumente und Einstellungen\jl.2G5\Desktop\C4D 8.5, SketchAndToon\8500\030911 8.500\resource\_api\c4d_resource.cpp   u�  s�  �'�'�    acos                  �?pow     ��    .?AVtype_info@@  �            �    .       @�S�S�S�S�S�S�S�S�SH    I�?          fmod         ������t�������������������0�0�0�0�0�0               ���5�h!����?      �?             ��       ���ܧ׹�fq�@      ��@�6C����?      �?exp          A�}�����          @T                            pT            �T            XT                                                                                                                        �            ������̙���[    �[                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �����������   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��  ���� 
                                     ��   X�	   ,�
   �   ܛ   ��   ��   \�   $�   ��   Ě   ��   d�x   T�y   D�z   4��   0��    �   ��   ��   ��   ��   ��   ��!   ��   ��   ��   |�   t�   l�   h�   d�    `�   X�   P�   H�   @�   8�   0�   (�    �   �"   �#   �$   �      �      ���������              �       �D        � 0         
      p?  �?   _       
          �?      �C      �;      �?      �?      ���tz�����������
.NSmr������6Jbv������:?Y^~������"6Nb�������     .      f5f5                    ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                ���5      @   �  �   ����                       �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �             x   
                                            	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �                       �  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��            �&  C   C                                                                                                                                   C                                                                                                                                   ��    �j���:�j|��:�hp��:Dfd��:od\��: _        
  040a    L�ESP D�ESP 850     1252      040b    <�FIN 4�FIN 850     1252      040c    ,�FRA $�FRA 850     1252      040f    �ISL �ISL 850     1252      041d    �SVE  �SWE 850     1252    -  042d    ��EUQ D�ESP 850     1252    
  080a    �ESM �MEX 850     1252      080c    ,�FRB ��BEL 850     1252      0c07    ؟DEA ПAUT 850     1252    	  0c09    ȟENA ��AUS 850     1252    
  0c0a    ��ESN D�ESP 850     1252      0c0c    ,�FRC ��CAN 850     1252    
  100a    �ESG ��GTM 850     1252      100c    ,�FRS ��CHE 850     1252    
  140a    �ESC x�CRI 850     1252      140c    ,�FRL l�LUX 850     1252    
  180a    �ESA d�PAN 850     1252    	  1c09    ȟENS T�ZAF 437     1252    
  1c0a    �ESD @�DOM 850     1252    
   200a    �ESV 4�VEN 850     1252    
$  240a    �ESO (�COL 850     1252    
(  280a    �ESR  �PER 850     1252    
,  2c0a    �ESS �ARG 850     1252    
0  300a    �ESF �ECU 850     1252    
4  340a    �ESL �CHL 850     1252    
8  380a    �ESY ��URY 850     1252    
<  3c0a    �ESZ �PRY 850     1252    6-T�USA L�GBR D�CHN <�CZE 4�GBR $�GBR �NLD �HKG �NZL  �NZL ��CHN �CHN ܠPRI ԠSVK ĠZAF ��KOR ��ZAF ��KOR ��TTO d�GBR x�GBR h�USA `�USA d�ENU P�ENU <�ENU 0�ENA (�NLB �ENC �ZHH �ZHI �CHS ��ZHH �CHS ФZHI ��CHT ��NLB ��ENU ��ENA |�ENL p�ENC \�ENB P�ENI @�ENJ 4�ENZ �ENS  �ENT ��ENG �ENU ܣENU ̣FRB ��FRC ��FRL ��FRS ��DEA t�DEC `�DEL P�DES @�ENI 0�ITS $�NOR �NOR ��NON �PTB ТESS ��ESB ��ESL ��ESO ��ESC l�ESD \�ESF H�ESE 4�ESG  �ESH �ESM  �ESN �ESI ܡESA ȡESZ ��ESR ��ESU ��ESY ��ESV p�SVF h�DES d�ENG `�ENU \�ENU �C    ��������������x�p�h�\�P�H�<�8�4�0�,�(�$� �����������(��إХĥ��������������x�             �@         �@         �@        @�@        P�@        $�@       ���@        ��@     ���4@   ������N@ �p+��ŝi@�]�%��O�@q�וC�)��@���D�����@�<զ��Ix��@o�����G���A��kU'9��p�|B�ݎ�����~�QC��v���)/��&D(�������D������Jz��Ee�Ǒ����Feu��uv�HMXB䧓9;5���SM��]=�];���Z�]�� �T��7a���Z��%]���g����'���]݀nLɛ� �R`�%u    �����������?q=
ףp=
ף�?Zd;�O��n��?��,e�X���?�#�GG�ŧ�?@��il��7��?3=�Bz�Ք���?����a�w̫�?/L[�Mľ����?��S;uD����?�g��9E��ϔ?$#�⼺;1a�z?aUY�~�S|�_?��/�����D?$?��9�'��*?}���d|F��U>c{�#Tw����=��:zc%C1��<!��8�G�� ��;܈X��ㆦ;ƄEB��u7�.:3q�#�2�I�Z9����Wڥ����2�h��R�DY�,%I�-64OS��k%�Y����}�����ZW�<�P�"NKeb�����}�-ޟ���ݦ�
�p     ����PST                                                             PDT                                                             �F8G����            ����            ����   ;   Z   x   �   �   �   �     0  N  m  ����   :   Y   w   �   �   �   �     /  M  l         ��    .?AVruntime_error@std@@ ��    .?AVfailure@ios_base@std@@      ��    .?AVios_base@std@@      ��    .?AVlogic_error@std@@   ��    .?AVlength_error@std@@  ��    .?AVout_of_range@std@@  ��    .?AVfacet@locale@std@@  ��    .?AV_Locimp@locale@std@@        ��    .?AV?$num_put@DV?$ostreambuf_iterator@DU?$char_traits@D@std@@@std@@@std@@       ��    .?AV?$numpunct@D@std@@                �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           h   ,1E13b3�3'4�4�4k5�5�56r6�678�8�8�8i9�9:�:�:�:�:j;�;�;�;�;<)<N<o<�<�<�<�<=�=�=>T>�>1?�?�?    T   a0�0F1�1
2�2%6f6�677p7z7�7�7�7�78%8�8�8�8�8�8�88:P:o:[;s;�;�;A<q<�<F=a=�= 0  8   X6C7�;�;�;�;9<X<a<z<�<=*=h=�>�>�>�>�>�>l?q?�?�? @  t   �0�0�0�0�0�0�0�0�0 1=2[2�23?4_4L56�7�89#9�9�:G;^;u;�;�;�;�;3<^<r<<�<==,=7===J=e=�=�=b>�>�>�>�>?.?�?   P  �   g0l0�0�0�0�0�0�0�0�0$1Y12B2t2�2�2�2�2�2�233333�3�3�3�3�34D4^4h4�4�4�4�4�4�4�4N5l5r5x5~5�5�5�566%6+616;6�6�6�6�6�6%7D7J7P7V7\7f7�7�8D9Q9�9�9�9�9�9:$:5:I:U:^=q==�=�>�>�>�?�?   `  0   �0�01E1]3{3�3�35�5�5�7�:�:;T;�;�<�>   p  t   K0g0�012A2[2u2�2�23�3I456@6s6�6�67?7r7�7�78>8q8�8�8
9=9p9�9�9	:b:P<a<r<�<�<�<�<�<F=N=`=r=�=>�>?2?M?�? �  x   0]0�0�01(1d1p1�1�1�1�12H2�2�2�23�3�3�3�34b4&5.5@5R5d5�5]6�6�627&8}8�8�8�97:J:O:b:~:�:�:�:;	;t;l=u=�=�=�=�= �  H   �1�1�1�2�2�2 3353g3�3�34$4,4Z4�4G5U5g5�8�86:�:&<(>�>�>0?^?�?�? �  D   ;0f0�0�1�1�1F23H3�3N5|5�5�5�5P7�7'858>9l9�9�9�9@;�;<%<Q?X? �  d   %3,3�3�5y7�7�7�7�7�78W8�8�8�8�899#9�;�;<+<|<�<=4=e=�=�=�=>d>�>�>�>�>�>�>?!?1?�?�?�?�? �  �   0/0L0x0�0�1�1�1�12(2H2�23T3k3{3�3<4S4c4�4)5@5P5l6�6�6�67S7q7�7�7*8�8�8�89*9T9v9�9�9::`:�:�:�:;;];�;�;h=�=�=�=>6>;>>l?�?   �  8   !0Q0w0�0�0!1�2�4�4�45S5�5�5�5�5�529h9f=�=�>�?�? �  0   E0n022�2�2�2�23`3�3�3@4�71;6;�;9=C=   �  L   �1�1�1�1�1N2z2�2�2�233N3�3�3T4�4�4�4�4 5�5�5�5�5�5�5E6�8�8�8�=�=     h   x2+3k3B4B:P:a:�:�:�:�:�:;�;�;�;�;�;�;<D<I<�<�<�<�<�<�<==&=x=�=�=�=�=�=�=>>X>t>�>�>H?\?�?�?  �   030@0P0n0v0�0�0�0�0�0�0,1O1�1�1�122,2t2�23%3.393L3U3q3y3�3�3�3�3+4�465�5788"8.848R8Z8�8�8�89�9�9�9	:�:�:�:;;';:;J;S;h;v;�;�;�;�;<G<_<�<�<�<�<�<�<�<�<�=�=�=�=1>�>�>?@?r?�?�?�?�?�?     �   00&010x0�0�0�0W1�1�1�1�1�12!2H2M2U2b2x2�23&3M3S3x3�3�3{4�4�4�4�4�4�4�455'5G5N5_5�5�5�5�56.6M6V6~6�6�6l7{7�7�7�7�7�7�7=8~8�8 939W9d9�9�9::P:�:�:�;�;r<�<=H=�=�==>�>�>�>?=?z?�?�?   0 �  �0�0\1�1�1'2f2�2�3�3�3�3�3�3�3�34464;4C4J4Q4j4q4x4�4�4�4�4�4�4�4�4�4�4�4�455!5(5=5F5N5V5^5f5n5v5~5�5�5�5�5�5�5�5�5�5�566�6�6�6�6�6 7\7�7�7888*838>8G8R8[8f8o8z8�8�8�8�8�8�8�8�8�8�8�8�8�8999#9.979B9K9V9_9j9s9~9�9�9�9�9�9�9�9�9�9�9�9�9�9
:::':2:;:F:O:Z:c:n:w:�:�:�:�:�:�:�:�: ;	;;;,;h;�;�;�;�;�;<<<"<+<6<?<J<S<^<g<v<�<�<*=f=�=�=�=�=�=�=>>>%>4>q>v>>�>�>�>�>�>�>�>�>�>�>�>�>????*?3?>?G?R?[?f?o?z?�?�?�?�?�?�?�?�?�?�?�?�?�? @   000#0.070B0K0V0_0j0s0~0�0�0�0�0�0�0�0�0�0�0�0�0�0
111'121;1F1O1Z1c1n1w1�1�1�1�1�1�1�1�1�1�1�1�1�1222"2+262?2J2S2^2g2r2{2�2�2�2�2�2�2�2�2�2�2�2�2�2333&3/3:3C3R3�3�3�3�3�3�3�3�3�3�3�3�3444 4)444=4H4Q4\4e4p4y4�4�4�4�4�4�4�4�4�45P5�5�5�5�5�5�5�5�50666=6L6�6�6�6�6�6�6�6.7g7l7u7�7�7�7�7�7�7�7�7�7888&8/8>8z8�8�8�8�8�8�8�8�8�899 9Y9^9g9r9{9�9�9::::%:0:9:D:M:X:a:l:u:�:�:�:�:�:�:�:�:�:�:�:�:�:;;; ;);4;=;H;Q;`;�;�;<L<R<Y<h<�<�<=X=�=�=>I>N>W>b>k>v>>�>�>�>�>�>�>�>????[?`?i?t?}?�?�?�?�?�?�?�?�?�?�?�?�? P    0	00Q0V0_0j0s0~0�0�0�01J1�1�1�1 2	222(212<2E2P2Y2h2�2�2�2�2�2�2�2�2�2�2333"3+3:3v3�3�3�3�3444%40494D4M4X4a4p4�4�4�4�4�4�4�4�4�45555*535>5G5R5[5f5o5z5�5�5�5�5�5�5�5�5�5�5�5�5�5666#6.676B6K6V6_6j6s6~6�6�6�6�6�6�6�6�6�6�6�6�6�6
777'727;7F7O7Z7c7n7w7�7�7�7�7�7�7�7�7�7�7�7�7�7888"8+868?8N8�8�89999%90999D9M9X9a9l9u9�9�9�9�9:::&:/:>:w:|:�:�:�:�:�:�:�:�:;;O;T;];h;q;|;�;�;�;�;�;�;�;�;�;�;�;�;�;<<<%<0<9<D<M<\<�<�<�<�<�<�<�<===V=�=�=
>F>�>�>�>�>???$?-?8?A?P?�?�?�?�?�?�?�?�? ` �  
000'020;0F0O0Z0c0n0w0�0�0�0�0�0�0�0�0�0�0�0�0�0111"1+161?1J1S1^1g1r1{1�1�1�1�1�1�1�1�1�1�1�1�1�1222&2/2:2C2N2W2b2k2v22�2�2�2�2�2�2�2�2�2�2�2�23333*333>3G3R3[3f3o3z3�3�3�3�3�3�3�3�3�3�3�3�3�3444#4.474B4K4V4_4j4s4~4�4�4�4�4�4�4�465r5�5�5&6_6d6m6x6�6�6�6�6�6�6�6�6�67E7J7S7^7g7r7{7�7�7�7�7�7�7�7�7888!808i8n8w8~8�8�8�8�8�8�8�8�859:9C9J9Q9X9�9�9:3:F:P:X:d:�:�:�:�:�: ;;#;K;�;�;�;�;&<?<R<�<=U=\=r=�=�=�=�=�=	>C>J>\>n>�>"?(?.?4?:?@?Q?a?�?�?�? p �   0A0Q0q0�0�0�0�0151Q1f1�1�1�1�1�1252T2�2�23j3�3b4�4�4�4�4515Q5q5�5�5�56!616Q6q6�6�6�6�6�6 7�7�78Q8}8�8�8�8919Q9q9�9�:;:;�;�;�;�;�;�;P<�<=A=Q=�=
>>>>:>Q>a>�>�>�>�>�>??1?]?�?�? � t   !0P0�0�0�0!1}1�12W24
44Z4b4�4�4�45J5�5�5�5�78H8�8�89Y9a9�9�9-:4:Q:q:�:�:�:;1;d;�;�;<M=�>�>q?�?�?�?�? � �   0�0�0�0�0�0�0c1�1�1E2a2q2�2�23�3�3�3�35!5A5a5}5�56:67�8�8�8�8�89"9I9�9 :b:�:�:�:�:�:;;*<4<><H<R<\<f<p<z<�<�<�=�=�=�=�=�=�=�=�=�=�=�=�=�=�>�>�>�>?(?a?�? � �   �1�1�123333#3*313e4�4�4�4�4�45<5@5D5H5L5P5a5q5�5�56)6/63686>6B6H6L6R6V6[6�6�637>7P7�7�7�7	8�8G9e9�9�9�9�9�9�9�9%:K:e:l:p:t:x:|:�:�:�:�:�:�:�:�:J;U;p;w;|;�;�;�;�;�;<<<<<<< <j<p<t<x<|<�<(=n=�=�=&>�> ?O?   � �   �01n1�1�1�1�13#3.353P3f3l3q3}3�3�3�3�3�3�5�5"6�6�6�6�6*7b7�7�7'8-8A8�889>9y99�9�9�9�9:::&:+:t:�:�:�:�:�:�:�:�:�:�:�:;;=;};�;�;�;�;E<�<�<>">1>9>D>J>P>Z>r>w>�>�>�>�>�>�>?h?�?�?�?�? � �   #0�0�0�0�0�0 111"1)1R1m1}1�1�1�2�24�5 6�67�7�8�8�899&9d9�9�9!:X:u:�:�:�:A;p;~;�;�;�;�;�;�;<#<;<K<�<>>D>L>T>\>h>m>y>�>�>�>�>�>�>�>�>�>�>?*?:?@?   � t   /343^4c4�5�5g7l7D8L8f8l8}8�8�8�8�8�8�8�8�8�899)9B9�9�9�9�9�9/:4:S:�:�:�:�:�:�:�:5;=;�;�;G<V<l<�=V>`?�?�?�? � �   T03 3$3(3,303438344)4�4�4�455*555I5O5]5f5w5�5�5�5�5�5�566+6N6Z6m6�6�6788$8f8x899x9�9:
:R:\:";,;�; <<<<<<E<k<�<�<�<�<�<�<�<�<�<�<�<�< ==j=u=�=�=�=�=�=�=�=>$>(>,>0>4>8><>@>�>�>�>�>�>�>   � �   ;0g0s0�0�0�0�0�0�0�0�0)1k1�1�1�1 2�2�2�2�2�2�2 3333;3G3O3W3g3~3�3�3�3�3�3�3�3�3�3�3�3�386F6L6f6k6z6�6�6�6�6�6�6�6�6�6�67777%7*7:7@7�7*8:":*:=:C:Y:`:f:p:v:{:�:�:�:�:�:�:�:@;�>�>�>??H?R?Z?`?h?q?z?   �    00003090C0I0c0i0q0�0�0�0%1?1�1�1�1�2�2�23h3�3�6�6�6�6�6�6�7�7�7�7�7�78>8H8i8~8�8�8�8999?9d9s9�9�9�9:::1:?:L:Q:W:�:�:;F;)<B<w<<�<�<�<�<D=W=�=�=�=�=�=�=	>>'>N>]>�>�>�>�>�>?$?+?7?�?    T   52_3e33�3�3�3�3�3�3�34[4�5�5�5�6�6�7�7�7�718�8+9;9G9Y9i9u9x:�:�:�:�:H;p;     @   u2�3�3%4�4�4�4-5q6�6�6�7�7�7U9d9�9�9�9�9�9+:c:u:�:�:W>m> 0 �   �12A2]2u2�2�2�2�2,3u3{3�3�3�3h4u4�4�4�4=5�5*6B6W6�6�6 777 7(7s7�7�7�7�8�8�89	99"9E9R9w9�9:%:2:o:�:�:�:�:;3;a;p;�;�;�;�;-<4<Z<r<�<�<�<�<�<�<p=k>�>�>??>? @ 0  /0G0�011.1l2�2�2�2�2�2�2�233>3D3e3o3z33�3�3�3�3�3�3�3444#4-474=4�4�4�4�4�4�4�4'5-5K5\5o5�5�5�5�5�5�5�566)6:6H6Q6W6c6h6r6y6�6�6�6�6�6�68888!8&8K8P8�8�8�8�8V9�9�9�9�9�9�9�9�9	::4:T:�:�: ;;;7;s;�;�;�;;<�<�<�<�<=t==�=�=�=�=�=�=�=>>.>8>S>\>a>h>p>z>�>�>�>�>�>�>�>�>A?S?�?�?�?�?�?   P �   w0191R1W1v1�1�1�1�1�1�1�1�12-2�2�2�263[3�5�56\6{6�6�6�67J7f778O8�8�8�9�9�9�9�9�9�9�9�9::	:�:�:�:;=�=�=�=�=�=�=:>l>�>�>�>?@?F?Q?]?f?l?p?{?�?�?�? ` P  t4}4�4�4�4�4�4�4�4�4�4 555!5.5?5D5K5Q5Y5_5g5q5v5�5�5�5�5�5�5�5�5�5�5�566'616:6F6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�677u8�8�8�8�8j9p9�9:X:`:e:x:}:�:�:�:�:�:�:�:�:?;Q;V;^;b;t;};�;�;�;�;�;�;�;�; <0<6<I<S<q<w<�<�<==)=<=D=K=S=_=j=q=w=|=�=�=�=�=�=>>0>8>>>F>N>]>o>u>|>�>�>�>�>�>�>�>�>�>???$?/?>?E?T?s?z?�?�?�?�?�?�?�?�?�?�?�?   p �   	00(070H0T0\0k0�0�0�0�0�0�0�0�0�0�0�011+1G1N1T1Y1m1u1z11�1�1�1�1�1�1%2E2P2�2�2�23!3,363@3J3T3	66�67�7�7�7	88!8=8P8W8i8q8�8�8�8�849z9�9~:�:�:�:);Y;�;�;�;&<K<f<�<�<�<�<�<=='=>=R=c=�=�=�=�=>>*>:>Q>i>z>�>�>a?�?�?�?�?�?�? � 0  090L0h0�0�0�0�01,1A1S1�1�1�1�1�1�1[2y2�2�2t3�3�3�3�3�3�3�3�3�3�3�3�3�3�34
4444%4C4l4t44�4�4�4�4 55Y5�5�5�5�5696D6b6�6�6�6�6�6!7-767B7K7V7b7}7�7�7�78$8>8o8t8~8�8�8�8�8�8�8�8�8�8989S9|9�9�9�9�9E:V:_:k:t::�:�:';P;v;�;�;�;�;�;�;<<<)<2<=<J<!=1=A=U=i=}=�=�=�=�=�=�=>!>5>I>g>y>�>�>�>?   � �  �2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2 33333333 3$3(3,3034383<3@3D3H3L3P3T3X3\3`3d3h3l3p3t3x3|3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3 44444444 4$4(4,404P4T4X4\4`4d4h4l4p4t4x4|4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4 55555555 5$5(5,5054585<5@5D5H5L5P5T5X5\5`5d5h5l5p5t5x5|5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5 66666666 6$6(6,6064686h6l6p6t6x6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6 77777777 7$7(7,7074787<7@7D7H7L7P7T7X7\7`7d7h7l7p7t7x7|7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7 8,888D8P8\8�8�8 99999$9(989@9D9P9X9\9�9�9�=>T>X>�>�>�>�>   � �  �6�6�6�6�6 777 7$7(7,7d7h7l7p7t7x7|7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7 88888888 8$8(8,80848@8X8l8|8�8�8�8�8�8�8�8�8 9999,90989<9T9d9h9p9�9�9�9�9�9�9�9�9�9::: :$:<:L:P:X:p:t:x:�:�:�:�:�:�:�:�:�:;;$;4;8;@;X;\;t;�;�;�;�;�;�;�;�;�;�;�;<$<(<4<H<T<h<t<x<�<�<�<�<�<�<�<�<(=<=H=P=�=�=�=�=�=�=�=�=�=�=�= >>(>D>L>P>\>d>p>�>�>�>�>�>�>?? ?,?@?L?P?T?\?d?p?�?�?�?�?�?�?�?�?�? � P   0$000L0T0h0t0x0|0�0�0�0�0�0�0�011141@1\1h1�1�1�1�1�1�1�1�1�1�122   � (   0000000 0$0(04080<0@0L0X0 �    �6�6   t   �<�<�<=8=H=L=P=T=X=\=`=d=h=l=x=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=z>~>�>�>�>�>�>�>P?d?h?l?p?x?       �1�1 22 0 h  2L2T2\2d2l2t2|2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�23333$3,343<3D3L3T3\3d3l3t3|3�3�3�3�3�3�3N4R4V4Z4^4b4f4j4n4r4v4z4~4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�455
555555"5&5*5.52565:5>5B5F5J5\5`5�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;<<8<@<d<l<�<�<�<�<�<�<==@=H=l=t=�=�=�=�=�=�=>$>H>P>t>|>�>�>�>�>�> ?$?,?P?X?|?�?�?�?�?�?   @ 8   00,040X0`0�0�0�0�0�0�0�0�0�0�0�0 1111 1(10181@1H1P1X1`1h1p1x1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 2222 2(20282@2H2P2X2`2h2p2x2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2 3333 3(30383@3H3P3X3`3h3p3x3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3 44444444 4$4(4x7|7808X8x8�8�8�8�8 9x9                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        